magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< pwell >>
rect 7068 22 7172 108
<< mvpsubdiff >>
rect 7094 48 7146 82
<< mvnsubdiff >>
rect 7119 1032 7171 1066
<< locali >>
rect 5546 2684 5580 2730
rect 5546 2604 5580 2650
rect 5546 2523 5580 2570
rect 5546 2442 5580 2489
rect 5546 2361 5580 2408
rect 5546 2280 5580 2327
rect 5702 2684 5736 2730
rect 5702 2604 5736 2650
rect 5702 2523 5736 2570
rect 5702 2442 5736 2489
rect 5702 2361 5736 2408
rect 5702 2280 5736 2327
rect 5622 2156 5660 2190
rect 24365 1237 24399 1275
rect 9768 1197 9809 1231
rect 9843 1197 9884 1231
rect 9918 1197 9959 1231
rect 9993 1197 10034 1231
rect 10068 1197 10109 1231
rect 10143 1197 10184 1231
rect 10218 1197 10259 1231
rect 10293 1197 10334 1231
rect 10368 1197 10409 1231
rect 10443 1197 10484 1231
rect 10518 1197 10559 1231
rect 10593 1197 10634 1231
rect 10668 1197 10709 1231
rect 10743 1197 10784 1231
rect 10818 1197 10858 1231
rect 10892 1197 10932 1231
rect 10966 1197 11006 1231
rect 11040 1197 11080 1231
rect 11114 1197 11154 1231
rect 11188 1197 11228 1231
<< viali >>
rect 5546 2730 5580 2764
rect 5546 2650 5580 2684
rect 5546 2570 5580 2604
rect 5546 2489 5580 2523
rect 5546 2408 5580 2442
rect 5546 2327 5580 2361
rect 5546 2246 5580 2280
rect 5702 2730 5736 2764
rect 5702 2650 5736 2684
rect 5702 2570 5736 2604
rect 5702 2489 5736 2523
rect 5702 2408 5736 2442
rect 5702 2327 5736 2361
rect 5702 2246 5736 2280
rect 5588 2156 5622 2190
rect 5660 2156 5694 2190
rect 24365 1275 24399 1309
rect 9734 1197 9768 1231
rect 9809 1197 9843 1231
rect 9884 1197 9918 1231
rect 9959 1197 9993 1231
rect 10034 1197 10068 1231
rect 10109 1197 10143 1231
rect 10184 1197 10218 1231
rect 10259 1197 10293 1231
rect 10334 1197 10368 1231
rect 10409 1197 10443 1231
rect 10484 1197 10518 1231
rect 10559 1197 10593 1231
rect 10634 1197 10668 1231
rect 10709 1197 10743 1231
rect 10784 1197 10818 1231
rect 10858 1197 10892 1231
rect 10932 1197 10966 1231
rect 11006 1197 11040 1231
rect 11080 1197 11114 1231
rect 11154 1197 11188 1231
rect 11228 1197 11262 1231
rect 24365 1203 24399 1237
<< metal1 >>
rect 5540 2764 5586 2776
rect 5540 2730 5546 2764
rect 5580 2730 5586 2764
rect 5540 2684 5586 2730
rect 5540 2650 5546 2684
rect 5580 2650 5586 2684
rect 5540 2604 5586 2650
rect 5540 2570 5546 2604
rect 5580 2570 5586 2604
rect 5540 2523 5586 2570
rect 5540 2489 5546 2523
rect 5580 2489 5586 2523
rect 5540 2442 5586 2489
rect 5540 2408 5546 2442
rect 5580 2408 5586 2442
rect 5540 2361 5586 2408
rect 5540 2327 5546 2361
rect 5580 2327 5586 2361
rect 5540 2280 5586 2327
rect 5540 2246 5546 2280
rect 5580 2246 5586 2280
rect 5540 2234 5586 2246
rect 5696 2764 5805 2776
rect 5696 2730 5702 2764
rect 5736 2730 5805 2764
rect 5696 2684 5805 2730
rect 5696 2650 5702 2684
rect 5736 2650 5805 2684
rect 5696 2604 5805 2650
rect 5696 2570 5702 2604
rect 5736 2570 5805 2604
rect 5696 2523 5805 2570
rect 5696 2489 5702 2523
rect 5736 2489 5805 2523
rect 5696 2442 5805 2489
rect 5696 2408 5702 2442
rect 5736 2408 5805 2442
rect 5696 2361 5805 2408
rect 5696 2327 5702 2361
rect 5736 2327 5805 2361
rect 5696 2280 5805 2327
rect 5696 2246 5702 2280
rect 5736 2246 5805 2280
rect 5696 2234 5805 2246
tri 5742 2214 5762 2234 ne
rect 5576 2190 5590 2196
rect 5576 2156 5588 2190
rect 5576 2150 5590 2156
rect 5584 2144 5590 2150
rect 5642 2144 5654 2196
rect 5706 2144 5712 2196
rect 4578 1922 4584 1974
rect 4636 1922 4648 1974
rect 4700 1922 5244 1974
tri 5202 1916 5208 1922 ne
rect 5208 1916 5244 1922
tri 5244 1916 5302 1974 sw
tri 5208 1895 5229 1916 ne
rect 4860 1881 4988 1887
rect 4860 1765 4868 1881
rect 4984 1765 4988 1881
rect 3542 1641 3707 1757
rect 3823 1641 3829 1757
rect 3542 1607 3637 1641
tri 3637 1607 3671 1641 nw
rect 2206 1298 2212 1350
rect 2264 1298 2276 1350
rect 2328 1298 2334 1350
tri 3522 1177 3542 1197 se
rect 3542 1177 3629 1607
tri 3629 1599 3637 1607 nw
rect 4609 1205 4779 1607
rect 4860 1329 4988 1765
rect 5030 1881 5082 1887
rect 5030 1817 5082 1829
rect 5030 1489 5082 1765
tri 5228 1573 5229 1574 se
rect 5229 1573 5302 1916
tri 5206 1551 5228 1573 se
rect 5228 1569 5302 1573
tri 5302 1569 5306 1573 sw
rect 5228 1551 5306 1569
rect 5206 1541 5306 1551
tri 5306 1541 5334 1569 sw
tri 5082 1489 5088 1495 sw
rect 5206 1489 5212 1541
rect 5264 1489 5276 1541
rect 5328 1489 5334 1541
rect 5030 1461 5088 1489
tri 5088 1461 5116 1489 sw
rect 5030 1409 5147 1461
rect 5199 1409 5211 1461
rect 5263 1409 5269 1461
tri 4988 1329 5002 1343 sw
rect 5131 1329 5137 1381
rect 5189 1329 5201 1381
rect 5253 1329 5327 1381
rect 4860 1309 5002 1329
tri 5002 1309 5022 1329 sw
tri 5259 1309 5279 1329 ne
rect 5279 1309 5327 1329
rect 4860 1301 5022 1309
tri 5022 1301 5030 1309 sw
tri 5279 1305 5283 1309 ne
rect 4860 1249 5123 1301
rect 5175 1249 5187 1301
rect 5239 1249 5245 1301
tri 3501 1156 3522 1177 se
rect 3522 1156 3629 1177
tri 5262 1156 5283 1177 se
rect 5283 1156 5327 1309
tri 5560 1237 5584 1261 se
rect 5584 1237 5655 2144
tri 5655 2109 5690 2144 nw
tri 5755 1649 5762 1656 se
rect 5762 1649 5805 2234
rect 5915 1948 5921 2000
rect 5973 1948 5985 2000
rect 6037 1948 6043 2000
tri 5917 1914 5951 1948 ne
tri 5805 1649 5812 1656 sw
tri 5727 1621 5755 1649 se
rect 5755 1621 5812 1649
tri 5812 1621 5840 1649 sw
rect 5726 1569 5732 1621
rect 5784 1569 5796 1621
rect 5848 1569 5854 1621
tri 5655 1237 5679 1261 sw
tri 5554 1231 5560 1237 se
rect 5560 1231 5679 1237
tri 5679 1231 5685 1237 sw
tri 5544 1221 5554 1231 se
rect 5554 1221 5685 1231
tri 5685 1221 5695 1231 sw
rect 5544 1169 5550 1221
rect 5602 1169 5637 1221
rect 5689 1169 5695 1221
rect 3501 1104 3507 1156
rect 3559 1104 3571 1156
rect 3623 1104 3629 1156
rect 3687 1104 3693 1156
rect 3745 1104 3757 1156
rect 3809 1145 5327 1156
rect 3809 1104 5286 1145
tri 5286 1104 5327 1145 nw
rect 5951 1156 6003 1948
tri 6351 1190 6352 1191 se
rect 6352 1190 6404 1833
tri 6404 1799 6438 1833 nw
tri 7870 1799 7901 1830 ne
rect 7901 1799 7956 1830
tri 7901 1798 7902 1799 ne
rect 7902 1798 7956 1799
tri 7956 1798 7988 1830 nw
rect 6468 1729 6557 1781
tri 6003 1156 6037 1190 sw
tri 6317 1156 6351 1190 se
rect 6351 1156 6404 1190
tri 6404 1156 6438 1190 sw
rect 5951 1104 5957 1156
rect 6009 1104 6021 1156
rect 6073 1104 6079 1156
rect 6310 1104 6316 1156
rect 6368 1104 6380 1156
rect 6432 1104 6438 1156
rect 6468 1186 6520 1729
tri 6520 1695 6554 1729 nw
rect 7320 1249 7326 1301
rect 7378 1249 7390 1301
rect 7442 1249 7448 1301
tri 6520 1186 6524 1190 sw
rect 6468 1156 6524 1186
tri 6524 1156 6554 1186 sw
rect 7320 1156 7448 1249
tri 7872 1156 7902 1186 se
rect 7902 1156 7954 1798
tri 7954 1796 7956 1798 nw
rect 22820 1787 22872 1793
rect 22820 1707 22872 1735
tri 22786 1426 22820 1460 se
rect 22820 1426 22872 1655
rect 20887 1329 20893 1381
rect 20945 1329 20957 1381
rect 21009 1329 21015 1381
rect 22727 1374 22733 1426
rect 22785 1374 22813 1426
rect 22865 1374 22872 1426
rect 8428 1249 8434 1301
rect 8486 1249 8498 1301
rect 8550 1249 8556 1301
rect 9722 1249 9728 1301
rect 9780 1249 9793 1301
rect 9845 1249 9858 1301
rect 9910 1249 9923 1301
rect 9975 1249 9988 1301
rect 10040 1249 10053 1301
rect 10105 1249 10118 1301
rect 10170 1249 10183 1301
rect 10235 1249 10248 1301
rect 10300 1249 10313 1301
rect 10365 1249 10378 1301
rect 10430 1249 10443 1301
rect 10495 1249 10508 1301
rect 10560 1249 10573 1301
rect 10625 1249 10638 1301
rect 10690 1249 10703 1301
rect 10755 1249 10768 1301
rect 10820 1249 10832 1301
rect 10884 1249 10896 1301
rect 10948 1249 10960 1301
rect 11012 1249 11024 1301
rect 11076 1249 11088 1301
rect 11140 1249 11152 1301
rect 11204 1249 11216 1301
rect 11268 1249 11274 1301
rect 9722 1231 11274 1249
rect 20887 1242 21015 1329
rect 24359 1319 24405 1321
rect 24356 1313 24408 1319
tri 22006 1270 22011 1275 se
rect 22011 1270 24217 1275
tri 21015 1242 21043 1270 sw
tri 21978 1242 22006 1270 se
rect 22006 1242 24217 1270
rect 9722 1197 9734 1231
rect 9768 1197 9809 1231
rect 9843 1197 9884 1231
rect 9918 1197 9959 1231
rect 9993 1197 10034 1231
rect 10068 1197 10109 1231
rect 10143 1197 10184 1231
rect 10218 1197 10259 1231
rect 10293 1197 10334 1231
rect 10368 1197 10409 1231
rect 10443 1197 10484 1231
rect 10518 1197 10559 1231
rect 10593 1197 10634 1231
rect 10668 1197 10709 1231
rect 10743 1197 10784 1231
rect 10818 1197 10858 1231
rect 10892 1197 10932 1231
rect 10966 1197 11006 1231
rect 11040 1197 11080 1231
rect 11114 1197 11154 1231
rect 11188 1197 11228 1231
rect 11262 1197 11274 1231
rect 9722 1191 11274 1197
rect 12664 1190 12670 1242
rect 12722 1190 12734 1242
rect 12786 1190 12794 1242
rect 20887 1190 20893 1242
rect 20945 1190 20957 1242
rect 21009 1237 21043 1242
tri 21043 1237 21048 1242 sw
tri 21973 1237 21978 1242 se
rect 21978 1237 24217 1242
rect 21009 1236 21048 1237
tri 21048 1236 21049 1237 sw
tri 21972 1236 21973 1237 se
rect 21973 1236 24217 1237
rect 21009 1190 21015 1236
tri 21950 1214 21972 1236 se
rect 21972 1214 24217 1236
rect 21679 1196 24217 1214
rect 21679 1191 23129 1196
tri 23129 1191 23134 1196 nw
tri 24081 1191 24086 1196 ne
rect 24086 1191 24217 1196
rect 24356 1249 24408 1261
rect 24356 1191 24408 1197
rect 21679 1190 23128 1191
tri 23128 1190 23129 1191 nw
tri 24086 1190 24087 1191 ne
rect 24087 1190 24217 1191
rect 6468 1104 6474 1156
rect 6526 1104 6538 1156
rect 6590 1104 6596 1156
rect 7320 1104 7326 1156
rect 7378 1104 7390 1156
rect 7442 1104 7448 1156
rect 7672 1104 7678 1156
rect 7730 1104 7742 1156
rect 7794 1139 7954 1156
rect 7794 1127 7942 1139
tri 7942 1127 7954 1139 nw
rect 21679 1182 23120 1190
tri 23120 1182 23128 1190 nw
tri 24087 1182 24095 1190 ne
rect 24095 1182 24217 1190
rect 7794 1104 7919 1127
tri 7919 1104 7942 1127 nw
rect 21679 1118 23056 1182
tri 23056 1118 23120 1182 nw
tri 24095 1149 24128 1182 ne
rect 24128 1152 24217 1182
tri 24217 1152 24247 1182 sw
rect 24128 1118 24247 1152
tri 24247 1118 24281 1152 sw
tri 25139 1118 25173 1152 se
rect 25173 1118 25373 1416
rect 21679 1108 23046 1118
tri 23046 1108 23056 1118 nw
rect 141 1070 341 1076
rect 193 1018 215 1070
rect 267 1018 289 1070
rect 141 1001 341 1018
rect 193 949 215 1001
rect 267 949 289 1001
rect 141 931 341 949
rect 193 879 215 931
rect 267 879 289 931
rect 141 873 341 879
rect 7058 873 7268 1076
rect 6855 839 7678 845
rect 6907 793 7678 839
rect 7730 793 7742 845
rect 7794 793 7800 845
rect 6855 775 6907 787
rect 5649 713 5655 765
rect 5707 713 5719 765
rect 5771 713 5777 765
tri 6907 759 6941 793 nw
rect 6855 717 6907 723
rect 7320 583 7372 589
rect 2002 476 2054 482
rect 268 405 274 457
rect 326 405 338 457
rect 390 405 398 457
rect 503 405 509 457
rect 561 405 573 457
rect 625 405 633 457
rect 1250 405 1257 457
rect 1309 405 1321 457
rect 1373 405 1380 457
rect 1713 405 1721 457
rect 1773 405 1785 457
rect 1837 405 1843 457
rect 2002 412 2054 424
rect 1250 402 1380 405
rect 2002 354 2054 360
rect 2838 405 2890 465
rect 2838 341 2890 353
rect 3577 454 3629 464
rect 3577 390 3629 402
rect 3577 332 3629 338
rect 3687 456 3739 464
rect 3687 392 3739 404
rect 3866 398 3918 525
rect 7320 519 7372 531
rect 6468 455 6520 464
rect 3687 334 3739 340
rect 6468 391 6520 403
rect 2838 283 2890 289
rect 6468 281 6520 339
rect 6855 456 6907 464
rect 6855 392 6907 404
rect 6855 334 6907 340
rect 6960 440 7012 464
rect 6960 376 7012 388
rect 7320 330 7372 467
rect 6960 318 7012 324
rect 7058 38 7556 253
rect 21679 50 21856 1108
tri 21856 1024 21940 1108 nw
rect 24128 958 25373 1118
rect 24128 938 24246 958
tri 24246 938 24266 958 nw
rect 23211 932 23263 938
rect 24128 910 24218 938
tri 24218 910 24246 938 nw
rect 23211 852 23263 880
tri 23205 794 23211 800 se
rect 23211 794 23263 800
tri 23163 752 23205 794 se
rect 23205 752 23263 794
rect 23174 724 23263 752
rect 23174 700 23239 724
tri 23239 700 23263 724 nw
rect 24413 361 24497 533
rect 5674 -122 5680 -70
rect 5732 -122 5744 -70
rect 5796 -122 6389 -70
<< via1 >>
rect 5590 2190 5642 2196
rect 5590 2156 5622 2190
rect 5622 2156 5642 2190
rect 5590 2144 5642 2156
rect 5654 2190 5706 2196
rect 5654 2156 5660 2190
rect 5660 2156 5694 2190
rect 5694 2156 5706 2190
rect 5654 2144 5706 2156
rect 4584 1922 4636 1974
rect 4648 1922 4700 1974
rect 4868 1765 4984 1881
rect 3707 1641 3823 1757
rect 2212 1298 2264 1350
rect 2276 1298 2328 1350
rect 5030 1829 5082 1881
rect 5030 1765 5082 1817
rect 5212 1489 5264 1541
rect 5276 1489 5328 1541
rect 5147 1409 5199 1461
rect 5211 1409 5263 1461
rect 5137 1329 5189 1381
rect 5201 1329 5253 1381
rect 5123 1249 5175 1301
rect 5187 1249 5239 1301
rect 5921 1948 5973 2000
rect 5985 1948 6037 2000
rect 5732 1569 5784 1621
rect 5796 1569 5848 1621
rect 5550 1169 5602 1221
rect 5637 1169 5689 1221
rect 3507 1104 3559 1156
rect 3571 1104 3623 1156
rect 3693 1104 3745 1156
rect 3757 1104 3809 1156
rect 5957 1104 6009 1156
rect 6021 1104 6073 1156
rect 6316 1104 6368 1156
rect 6380 1104 6432 1156
rect 7326 1249 7378 1301
rect 7390 1249 7442 1301
rect 22820 1735 22872 1787
rect 22820 1655 22872 1707
rect 20893 1329 20945 1381
rect 20957 1329 21009 1381
rect 22733 1374 22785 1426
rect 22813 1374 22865 1426
rect 8434 1249 8486 1301
rect 8498 1249 8550 1301
rect 9728 1249 9780 1301
rect 9793 1249 9845 1301
rect 9858 1249 9910 1301
rect 9923 1249 9975 1301
rect 9988 1249 10040 1301
rect 10053 1249 10105 1301
rect 10118 1249 10170 1301
rect 10183 1249 10235 1301
rect 10248 1249 10300 1301
rect 10313 1249 10365 1301
rect 10378 1249 10430 1301
rect 10443 1249 10495 1301
rect 10508 1249 10560 1301
rect 10573 1249 10625 1301
rect 10638 1249 10690 1301
rect 10703 1249 10755 1301
rect 10768 1249 10820 1301
rect 10832 1249 10884 1301
rect 10896 1249 10948 1301
rect 10960 1249 11012 1301
rect 11024 1249 11076 1301
rect 11088 1249 11140 1301
rect 11152 1249 11204 1301
rect 11216 1249 11268 1301
rect 24356 1309 24408 1313
rect 24356 1275 24365 1309
rect 24365 1275 24399 1309
rect 24399 1275 24408 1309
rect 12670 1190 12722 1242
rect 12734 1190 12786 1242
rect 20893 1190 20945 1242
rect 20957 1190 21009 1242
rect 24356 1261 24408 1275
rect 24356 1237 24408 1249
rect 24356 1203 24365 1237
rect 24365 1203 24399 1237
rect 24399 1203 24408 1237
rect 24356 1197 24408 1203
rect 6474 1104 6526 1156
rect 6538 1104 6590 1156
rect 7326 1104 7378 1156
rect 7390 1104 7442 1156
rect 7678 1104 7730 1156
rect 7742 1104 7794 1156
rect 141 1018 193 1070
rect 215 1018 267 1070
rect 289 1018 341 1070
rect 141 949 193 1001
rect 215 949 267 1001
rect 289 949 341 1001
rect 141 879 193 931
rect 215 879 267 931
rect 289 879 341 931
rect 6855 787 6907 839
rect 7678 793 7730 845
rect 7742 793 7794 845
rect 5655 713 5707 765
rect 5719 713 5771 765
rect 6855 723 6907 775
rect 7320 531 7372 583
rect 274 405 326 457
rect 338 405 390 457
rect 509 405 561 457
rect 573 405 625 457
rect 1257 405 1309 457
rect 1321 405 1373 457
rect 1721 405 1773 457
rect 1785 405 1837 457
rect 2002 424 2054 476
rect 2002 360 2054 412
rect 2838 353 2890 405
rect 2838 289 2890 341
rect 3577 402 3629 454
rect 3577 338 3629 390
rect 3687 404 3739 456
rect 7320 467 7372 519
rect 6468 403 6520 455
rect 3687 340 3739 392
rect 6468 339 6520 391
rect 6855 404 6907 456
rect 6855 340 6907 392
rect 6960 388 7012 440
rect 6960 324 7012 376
rect 23211 880 23263 932
rect 23211 800 23263 852
rect 5680 -122 5732 -70
rect 5744 -122 5796 -70
<< metal2 >>
rect 88 3118 5739 3318
rect 8514 3139 9382 3297
rect 88 1249 288 3118
tri 288 2906 500 3118 nw
rect 9965 2913 10137 2997
rect 22664 2246 22784 2339
rect 5584 2144 5590 2196
rect 5642 2144 5654 2196
rect 5706 2144 5712 2196
tri 3535 1922 3587 1974 se
rect 3587 1922 4584 1974
rect 4636 1922 4648 1974
rect 4700 1922 4706 1974
rect 5915 1948 5921 2000
rect 5973 1948 5985 2000
rect 6037 1948 6043 2000
tri 3523 1910 3535 1922 se
rect 3535 1910 3613 1922
tri 3613 1910 3625 1922 nw
rect 3523 1881 3584 1910
tri 3584 1881 3613 1910 nw
tri 4854 1881 4860 1887 se
rect 4860 1881 4988 1887
rect 532 1383 648 1637
rect 532 1267 770 1383
tri 3505 1350 3523 1368 se
rect 3523 1352 3581 1881
tri 3581 1878 3584 1881 nw
tri 4851 1878 4854 1881 se
rect 4854 1878 4868 1881
tri 4823 1850 4851 1878 se
rect 4851 1850 4868 1878
rect 3701 1765 4868 1850
rect 4984 1765 4988 1881
rect 3701 1758 4988 1765
rect 5030 1881 5082 1887
rect 5030 1817 5082 1829
rect 5030 1759 5082 1765
rect 22820 1787 22872 1793
rect 3701 1757 3881 1758
tri 3881 1757 3882 1758 nw
rect 3701 1641 3707 1757
rect 3823 1735 3859 1757
tri 3859 1735 3881 1757 nw
rect 3823 1707 3831 1735
tri 3831 1707 3859 1735 nw
rect 22820 1707 22872 1735
rect 3823 1641 3829 1707
tri 3829 1705 3831 1707 nw
rect 22820 1649 22872 1655
rect 5726 1569 5732 1621
rect 5784 1569 5796 1621
rect 5848 1569 5854 1621
rect 5206 1489 5212 1541
rect 5264 1489 5276 1541
rect 5328 1489 5661 1541
tri 21938 1489 21942 1493 se
rect 21942 1489 23339 1493
tri 21913 1464 21938 1489 se
rect 21938 1464 23339 1489
tri 23339 1464 23368 1493 sw
tri 21910 1461 21913 1464 se
rect 21913 1463 23368 1464
rect 21913 1461 21942 1463
rect 5141 1409 5147 1461
rect 5199 1409 5211 1461
rect 5263 1409 5661 1461
tri 21889 1440 21910 1461 se
rect 21910 1440 21942 1461
tri 21942 1440 21965 1463 nw
tri 23316 1440 23339 1463 ne
rect 23339 1440 23368 1463
tri 21875 1426 21889 1440 se
rect 21889 1426 21928 1440
tri 21928 1426 21942 1440 nw
tri 23339 1426 23353 1440 ne
rect 23353 1426 23368 1440
tri 23368 1426 23406 1464 sw
tri 21858 1409 21875 1426 se
rect 21875 1409 21889 1426
tri 21836 1387 21858 1409 se
rect 21858 1387 21889 1409
tri 21889 1387 21928 1426 nw
tri 21830 1381 21836 1387 se
rect 21836 1381 21876 1387
rect 3523 1350 3579 1352
tri 3579 1350 3581 1352 nw
rect 2206 1298 2212 1350
rect 2264 1298 2276 1350
rect 2328 1329 3558 1350
tri 3558 1329 3579 1350 nw
rect 5131 1329 5137 1381
rect 5189 1329 5201 1381
rect 5253 1329 20893 1381
rect 20945 1329 20957 1381
rect 21009 1329 21052 1381
tri 21823 1374 21830 1381 se
rect 21830 1374 21876 1381
tri 21876 1374 21889 1387 nw
rect 22727 1374 22733 1426
rect 22785 1374 22813 1426
rect 22865 1398 23235 1426
tri 23235 1398 23263 1426 sw
tri 23353 1411 23368 1426 ne
rect 23368 1411 23406 1426
tri 23406 1411 23421 1426 sw
rect 22865 1374 23263 1398
tri 21783 1334 21823 1374 se
rect 21823 1334 21836 1374
tri 21836 1334 21876 1374 nw
tri 23164 1334 23204 1374 ne
rect 23204 1334 23263 1374
tri 23368 1358 23421 1411 ne
tri 23421 1358 23474 1411 sw
tri 21778 1329 21783 1334 se
rect 21783 1329 21829 1334
rect 2328 1327 3556 1329
tri 3556 1327 3558 1329 nw
tri 21776 1327 21778 1329 se
rect 21778 1327 21829 1329
tri 21829 1327 21836 1334 nw
tri 23204 1327 23211 1334 ne
rect 2328 1313 3542 1327
tri 3542 1313 3556 1327 nw
tri 21762 1313 21776 1327 se
rect 21776 1313 21815 1327
tri 21815 1313 21829 1327 nw
rect 2328 1301 3530 1313
tri 3530 1301 3542 1313 nw
tri 21750 1301 21762 1313 se
rect 21762 1301 21803 1313
tri 21803 1301 21815 1313 nw
rect 2328 1298 3527 1301
tri 3527 1298 3530 1301 nw
tri 288 1249 299 1260 sw
rect 5117 1249 5123 1301
rect 5175 1249 5187 1301
rect 5239 1249 7326 1301
rect 7378 1249 7390 1301
rect 7442 1249 7448 1301
rect 8428 1249 8434 1301
rect 8486 1249 8498 1301
rect 8550 1249 9728 1301
rect 9780 1249 9793 1301
rect 9845 1249 9858 1301
rect 9910 1249 9923 1301
rect 9975 1249 9988 1301
rect 10040 1249 10053 1301
rect 10105 1249 10118 1301
rect 10170 1249 10183 1301
rect 10235 1249 10248 1301
rect 10300 1249 10313 1301
rect 10365 1249 10378 1301
rect 10430 1249 10443 1301
rect 10495 1249 10508 1301
rect 10560 1249 10573 1301
rect 10625 1249 10638 1301
rect 10690 1249 10703 1301
rect 10755 1249 10768 1301
rect 10820 1249 10832 1301
rect 10884 1249 10896 1301
rect 10948 1249 10960 1301
rect 11012 1249 11024 1301
rect 11076 1249 11088 1301
rect 11140 1249 11152 1301
rect 11204 1249 11216 1301
rect 11268 1249 11274 1301
tri 12683 1261 12723 1301 se
rect 12723 1271 21773 1301
tri 21773 1271 21803 1301 nw
rect 12723 1261 12813 1271
tri 12813 1261 12823 1271 nw
tri 12671 1249 12683 1261 se
rect 12683 1249 12801 1261
tri 12801 1249 12813 1261 nw
rect 88 1242 299 1249
tri 299 1242 306 1249 sw
tri 12664 1242 12671 1249 se
rect 12671 1242 12794 1249
tri 12794 1242 12801 1249 nw
rect 88 1227 306 1242
tri 306 1227 321 1242 sw
tri 12649 1227 12664 1242 se
rect 12664 1227 12670 1242
rect 88 1221 321 1227
tri 321 1221 327 1227 sw
tri 11473 1221 11479 1227 se
rect 11479 1221 12670 1227
rect 88 1215 327 1221
tri 327 1215 333 1221 sw
rect 88 1169 333 1215
tri 333 1169 379 1215 sw
rect 2926 1184 5550 1221
rect 88 1156 379 1169
tri 379 1156 392 1169 sw
rect 88 1104 392 1156
tri 392 1104 444 1156 sw
tri 2910 1104 2926 1120 se
rect 2926 1104 2978 1184
tri 2978 1172 2990 1184 nw
tri 5528 1172 5540 1184 ne
rect 5540 1172 5550 1184
tri 5540 1169 5543 1172 ne
rect 5543 1169 5550 1172
rect 5602 1169 5637 1221
rect 5689 1190 12670 1221
rect 12722 1190 12734 1242
rect 12786 1190 12794 1242
rect 20887 1190 20893 1242
rect 20945 1190 20957 1242
rect 21009 1190 21015 1242
rect 5689 1184 11503 1190
tri 11503 1184 11509 1190 nw
rect 5689 1169 5695 1184
tri 5695 1169 5710 1184 nw
rect 3501 1104 3507 1156
rect 3559 1104 3571 1156
rect 3623 1104 3629 1156
rect 88 1076 444 1104
tri 444 1076 472 1104 sw
tri 2882 1076 2910 1104 se
rect 2910 1076 2978 1104
rect 88 1070 472 1076
tri 2029 1070 2035 1076 se
rect 2035 1070 2978 1076
tri 3543 1070 3577 1104 ne
rect 88 1018 141 1070
rect 193 1018 215 1070
rect 267 1018 289 1070
rect 341 1018 472 1070
rect 88 1001 472 1018
rect 88 949 141 1001
rect 193 949 215 1001
rect 267 949 289 1001
rect 341 949 472 1001
rect 88 931 472 949
rect 88 879 141 931
rect 193 879 215 931
rect 267 879 289 931
rect 341 879 472 931
rect 88 873 472 879
tri 2002 1043 2029 1070 se
rect 2029 1049 2978 1070
rect 2029 1043 2972 1049
tri 2972 1043 2978 1049 nw
rect 2002 1027 2956 1043
tri 2956 1027 2972 1043 nw
rect 2002 476 2054 1027
tri 2054 1004 2077 1027 nw
rect 148 405 274 457
rect 326 405 338 457
rect 390 405 396 457
rect 503 405 509 457
rect 561 405 573 457
rect 625 405 631 457
rect 1251 405 1257 457
rect 1309 405 1321 457
rect 1373 405 1667 457
rect 1715 405 1721 457
rect 1773 405 1785 457
rect 1837 405 1843 457
rect 148 398 246 405
tri 246 398 253 405 nw
rect 503 398 584 405
tri 584 398 591 405 nw
tri 1581 398 1588 405 ne
rect 1588 398 1667 405
rect 148 371 219 398
tri 219 371 246 398 nw
tri 476 371 503 398 se
rect 503 371 557 398
tri 557 371 584 398 nw
tri 1588 371 1615 398 ne
rect 148 360 208 371
tri 208 360 219 371 nw
tri 465 360 476 371 se
rect 476 360 546 371
tri 546 360 557 371 nw
rect 148 353 201 360
tri 201 353 208 360 nw
tri 458 353 465 360 se
rect 465 353 539 360
tri 539 353 546 360 nw
rect 148 -122 200 353
tri 200 352 201 353 nw
tri 457 352 458 353 se
rect 458 352 527 353
tri 446 341 457 352 se
rect 457 341 527 352
tri 527 341 539 353 nw
tri 422 317 446 341 se
rect 446 317 503 341
tri 503 317 527 341 nw
tri 394 289 422 317 se
rect 422 289 475 317
tri 475 289 503 317 nw
tri 383 278 394 289 se
rect 394 278 464 289
tri 464 278 475 289 nw
rect 383 38 435 278
tri 435 249 464 278 nw
rect 1615 49 1667 398
tri 1723 371 1757 405 ne
rect 1757 198 1809 405
tri 1809 371 1843 405 nw
rect 2002 412 2054 424
rect 3577 454 3629 1104
rect 2002 354 2054 360
rect 2838 405 2890 411
rect 2838 341 2890 353
rect 3577 390 3629 402
rect 3577 332 3629 338
rect 3687 1104 3693 1156
rect 3745 1104 3757 1156
rect 3809 1104 3815 1156
rect 4434 1140 5501 1156
tri 5501 1140 5517 1156 sw
tri 5742 1140 5758 1156 se
rect 5758 1140 5957 1156
rect 4434 1104 5957 1140
rect 6009 1104 6021 1156
rect 6073 1104 6079 1156
rect 6310 1104 6316 1156
rect 6368 1104 6380 1156
rect 6432 1104 6438 1156
rect 3687 456 3739 1104
tri 3739 1070 3773 1104 nw
rect 4434 1078 4495 1104
tri 4495 1078 4521 1104 nw
tri 4428 713 4434 719 se
rect 4434 713 4487 1078
tri 4487 1070 4495 1078 nw
tri 6302 1070 6310 1078 se
rect 6310 1070 6438 1104
tri 6282 1050 6302 1070 se
rect 6302 1050 6438 1070
tri 4400 685 4428 713 se
rect 4428 685 4487 713
rect 5362 1026 6438 1050
rect 5362 999 6411 1026
tri 6411 999 6438 1026 nw
rect 6468 1104 6474 1156
rect 6526 1104 6538 1156
rect 6590 1104 6596 1156
rect 7320 1104 7326 1156
rect 7378 1104 7390 1156
rect 7442 1104 7448 1156
rect 7672 1104 7678 1156
rect 7730 1104 7742 1156
rect 7794 1104 7800 1156
rect 5362 454 5414 999
tri 5414 965 5448 999 nw
rect 5649 713 5655 765
rect 5707 713 5719 765
rect 5771 713 5777 765
tri 5649 700 5662 713 ne
rect 5662 700 5743 713
tri 5743 700 5756 713 nw
rect 3687 392 3739 404
rect 3687 334 3739 340
rect 2890 289 5620 302
rect 2838 250 5620 289
rect 1757 146 5516 198
rect 1914 66 5412 118
tri 1667 49 1683 65 sw
rect 1615 44 1683 49
tri 1615 38 1621 44 ne
rect 1621 38 1683 44
tri 1683 38 1694 49 sw
rect 5360 40 5412 66
rect 5464 38 5516 146
rect 5568 38 5620 250
tri 1621 -24 1683 38 ne
rect 1683 -24 1694 38
tri 1694 -24 1756 38 sw
tri 1683 -40 1699 -24 ne
tri 1698 -127 1699 -126 se
rect 1699 -127 1756 -24
rect 5662 -70 5714 700
tri 5714 671 5743 700 nw
rect 5782 346 5834 474
tri 5748 339 5755 346 ne
rect 5755 339 5834 346
tri 5755 333 5761 339 ne
rect 5761 333 5834 339
rect 6468 455 6520 1104
tri 6520 1070 6554 1104 nw
rect 6468 391 6520 403
rect 6468 333 6520 339
rect 6855 839 6907 845
rect 6855 775 6907 787
rect 6855 456 6907 723
rect 7320 583 7372 1104
tri 7372 1070 7406 1104 nw
rect 7672 852 7724 1104
tri 7724 1070 7758 1104 nw
rect 23211 932 23263 1334
tri 23421 1313 23466 1358 ne
rect 23466 1319 23474 1358
tri 23474 1319 23513 1358 sw
rect 23466 1313 23513 1319
tri 23513 1313 23519 1319 sw
rect 24356 1313 24408 1319
tri 23466 1305 23474 1313 ne
rect 23474 1305 23519 1313
tri 23519 1305 23527 1313 sw
tri 23474 1261 23518 1305 ne
rect 23518 1283 23527 1305
tri 23527 1283 23549 1305 sw
rect 23518 1261 23549 1283
tri 23549 1261 23571 1283 sw
tri 24334 1261 24356 1283 se
tri 23518 1252 23527 1261 ne
rect 23527 1252 23571 1261
tri 23571 1252 23580 1261 sw
tri 24325 1252 24334 1261 se
rect 24334 1252 24408 1261
tri 23527 1249 23530 1252 ne
rect 23530 1249 24408 1252
tri 23530 1222 23557 1249 ne
rect 23557 1222 24356 1249
tri 24325 1197 24350 1222 ne
rect 24350 1197 24356 1222
tri 24350 1191 24356 1197 ne
rect 24356 1191 24408 1197
tri 7724 852 7751 879 sw
rect 23211 852 23263 880
rect 7672 845 7751 852
tri 7751 845 7758 852 sw
rect 7672 793 7678 845
rect 7730 793 7742 845
rect 7794 793 7800 845
rect 24253 835 24368 880
rect 23211 794 23263 800
rect 23870 646 23974 685
rect 7320 519 7372 531
rect 7320 461 7372 467
rect 6855 392 6907 404
rect 6855 334 6907 340
rect 6960 440 7012 446
rect 6960 376 7012 388
tri 5761 324 5770 333 ne
rect 5770 324 5834 333
tri 5770 312 5782 324 ne
rect 5782 10 5834 324
rect 6960 38 7012 324
rect 7836 169 7845 225
rect 7901 169 7929 225
rect 7985 169 8013 225
rect 8069 169 8098 225
rect 8154 169 8163 225
rect 7836 93 8163 169
rect 7836 37 7845 93
rect 7901 37 7929 93
rect 7985 37 8013 93
rect 8069 37 8098 93
rect 8154 37 8163 93
rect 13533 60 14080 198
tri 5714 -70 5748 -36 sw
rect 5674 -122 5680 -70
rect 5732 -122 5744 -70
rect 5796 -122 5802 -70
tri 1675 -150 1698 -127 se
rect 1698 -150 1756 -127
tri 1756 -150 1779 -127 sw
<< via2 >>
rect 7845 169 7901 225
rect 7929 169 7985 225
rect 8013 169 8069 225
rect 8098 169 8154 225
rect 7845 37 7901 93
rect 7929 37 7985 93
rect 8013 37 8069 93
rect 8098 37 8154 93
<< metal3 >>
rect 8757 3244 8831 3318
rect 9986 1082 10158 1166
rect 7833 225 8166 230
rect 7833 169 7845 225
rect 7901 169 7929 225
rect 7985 169 8013 225
rect 8069 169 8098 225
rect 8154 169 8166 225
rect 7833 93 8166 169
rect 7833 37 7845 93
rect 7901 37 7929 93
rect 7985 37 8013 93
rect 8069 37 8098 93
rect 8154 37 8166 93
tri 7485 -4092 7833 -3744 se
rect 7833 -3932 8166 37
rect 7833 -4092 8006 -3932
tri 8006 -4092 8166 -3932 nw
rect 7485 -5000 7873 -4092
tri 7873 -4225 8006 -4092 nw
use sky130_fd_io__gpio_ovtv2_buf_localesd  sky130_fd_io__gpio_ovtv2_buf_localesd_0
timestamp 1648127584
transform 0 -1 5443 -1 0 3318
box 0 0 2114 5443
use sky130_fd_io__gpio_ovtv2_ibuf_se  sky130_fd_io__gpio_ovtv2_ibuf_se_0
timestamp 1648127584
transform 1 0 5647 0 1 0
box -2286 -894 19746 3465
use sky130_fd_io__gpio_ovtv2_ictl_logic  sky130_fd_io__gpio_ovtv2_ictl_logic_0
timestamp 1648127584
transform 1 0 141 0 1 12
box 0 -134 7045 1121
<< labels >>
flabel metal3 s 9986 1082 10158 1166 3 FreeSans 200 0 0 0 VCCHIB
port 1 nsew
flabel metal3 s 8757 3244 8831 3318 3 FreeSans 520 90 0 0 ENABLE_VDDIO_LV
port 2 nsew
flabel metal3 s 10072 1124 10072 1124 3 FreeSans 200 0 0 0 VCCHIB
port 1 nsew
flabel metal1 s 24413 361 24497 533 3 FreeSans 200 90 0 0 VCCHIB
port 1 nsew
flabel metal1 s 4629 1273 4761 1477 3 FreeSans 200 0 0 0 PAD
port 3 nsew
flabel metal2 s 9965 2913 10137 2997 3 FreeSans 200 0 0 0 VCCHIB
port 1 nsew
flabel metal2 s 13533 60 14080 198 3 FreeSans 200 0 0 0 VSSD
port 4 nsew
flabel metal2 s 8514 3139 9382 3297 3 FreeSans 200 0 0 0 VDDIO_Q
port 5 nsew
flabel metal2 s 22664 2246 22784 2339 3 FreeSans 200 0 0 0 VINREF
port 6 nsew
flabel metal2 s 24253 835 24368 880 3 FreeSans 200 0 0 0 OUT_H
port 7 nsew
flabel metal2 s 23870 646 23974 685 3 FreeSans 200 0 0 0 OUT
port 8 nsew
flabel metal2 s 6960 38 7012 103 3 FreeSans 200 0 0 0 HYS_TRIM_H
port 9 nsew
flabel metal2 s 5662 38 5714 128 3 FreeSans 200 0 0 0 IB_MODE_SEL_H[1]
port 10 nsew
flabel metal2 s 5783 38 5834 124 3 FreeSans 200 0 0 0 IB_MODE_SEL_H[0]
port 11 nsew
flabel metal2 s 2838 318 2890 406 3 FreeSans 200 0 0 0 VTRIP_SEL_H
port 12 nsew
flabel metal2 s 1757 371 1809 439 3 FreeSans 200 0 0 0 INP_DIS_H_N
port 13 nsew
flabel metal2 s 1615 49 1667 115 3 FreeSans 200 0 0 0 DM_H_N[2]
port 14 nsew
flabel metal2 s 148 38 200 113 3 FreeSans 200 0 0 0 DM_H_N[1]
port 15 nsew
flabel metal2 s 383 38 435 104 3 FreeSans 200 0 0 0 DM_H_N[0]
port 16 nsew
<< properties >>
string GDS_END 36591476
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 36564056
<< end >>
