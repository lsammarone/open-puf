/farmshare/home/classes/ee/372/PDKs/share/pdk/sky130A/libs.ref/sky130_fd_io/spice/sky130_ef_io__analog_pad.spice