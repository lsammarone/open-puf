magic
tech sky130A
timestamp 1649788711
use sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p15  sky130_fd_pr__rf_nfet_01v8_aM02W1p65L0p15_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1648127584
transform 1 0 451 0 1 -498
box 5 5 257 262
use sky130_fd_pr__pfet_01v8_lvt_A7J7BP  xm1
timestamp 1649788711
transform 1 0 0 0 1 1000
box -147 -695 147 695
use sky130_fd_pr__nfet_01v8_lvt_3WARGN  xm2
timestamp 1649788711
transform 1 0 0 0 1 -1000
box -129 -494 129 494
<< end >>
