magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 275 157 459 203
rect 1 21 459 157
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 151 47 181 131
rect 223 47 253 131
rect 351 47 381 177
<< scpmoshvt >>
rect 79 300 109 384
rect 163 300 193 384
rect 256 300 286 384
rect 351 297 381 497
<< ndiff >>
rect 301 131 351 177
rect 27 93 79 131
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 47 151 131
rect 181 47 223 131
rect 253 109 351 131
rect 253 75 307 109
rect 341 75 351 109
rect 253 47 351 75
rect 381 119 433 177
rect 381 85 391 119
rect 425 85 433 119
rect 381 47 433 85
<< pdiff >>
rect 299 485 351 497
rect 299 451 307 485
rect 341 451 351 485
rect 299 438 351 451
rect 301 384 351 438
rect 27 346 79 384
rect 27 312 35 346
rect 69 312 79 346
rect 27 300 79 312
rect 109 376 163 384
rect 109 342 119 376
rect 153 342 163 376
rect 109 300 163 342
rect 193 357 256 384
rect 193 323 212 357
rect 246 323 256 357
rect 193 300 256 323
rect 286 300 351 384
rect 301 297 351 300
rect 381 471 433 497
rect 381 437 391 471
rect 425 437 433 471
rect 381 403 433 437
rect 381 369 391 403
rect 425 369 433 403
rect 381 297 433 369
<< ndiffc >>
rect 35 59 69 93
rect 307 75 341 109
rect 391 85 425 119
<< pdiffc >>
rect 307 451 341 485
rect 35 312 69 346
rect 119 342 153 376
rect 212 323 246 357
rect 391 437 425 471
rect 391 369 425 403
<< poly >>
rect 351 497 381 523
rect 163 476 217 492
rect 163 442 173 476
rect 207 442 217 476
rect 163 426 217 442
rect 79 384 109 425
rect 163 384 193 426
rect 256 384 286 410
rect 79 251 109 300
rect 163 282 193 300
rect 25 203 109 251
rect 25 169 35 203
rect 69 169 109 203
rect 25 146 109 169
rect 79 131 109 146
rect 151 257 193 282
rect 256 259 286 300
rect 351 265 381 297
rect 151 131 181 257
rect 235 243 289 259
rect 235 226 245 243
rect 223 209 245 226
rect 279 209 289 243
rect 223 193 289 209
rect 331 249 385 265
rect 331 215 341 249
rect 375 215 385 249
rect 331 199 385 215
rect 223 170 265 193
rect 351 177 381 199
rect 223 146 260 170
rect 223 131 253 146
rect 79 21 109 47
rect 151 21 181 47
rect 223 21 253 47
rect 351 21 381 47
<< polycont >>
rect 173 442 207 476
rect 35 169 69 203
rect 245 209 279 243
rect 341 215 375 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 17 416 138 527
rect 173 476 269 493
rect 207 442 269 476
rect 173 425 269 442
rect 303 485 354 527
rect 303 451 307 485
rect 341 451 354 485
rect 303 418 354 451
rect 388 471 443 493
rect 388 437 391 471
rect 425 437 443 471
rect 17 396 140 416
rect 103 391 140 396
rect 388 403 443 437
rect 103 376 169 391
rect 17 346 69 362
rect 17 312 35 346
rect 103 342 119 376
rect 153 342 169 376
rect 203 357 354 377
rect 203 327 212 357
rect 200 323 212 327
rect 246 323 354 357
rect 388 369 391 403
rect 425 369 443 403
rect 388 353 443 369
rect 200 320 354 323
rect 197 318 354 320
rect 196 315 375 318
rect 192 312 375 315
rect 17 272 69 312
rect 188 310 375 312
rect 183 308 375 310
rect 169 302 375 308
rect 165 296 375 302
rect 161 290 375 296
rect 155 285 375 290
rect 148 278 375 285
rect 142 277 375 278
rect 142 276 220 277
rect 142 274 215 276
rect 142 273 212 274
rect 142 272 209 273
rect 17 271 209 272
rect 17 269 207 271
rect 17 268 205 269
rect 17 266 203 268
rect 17 264 202 266
rect 17 263 201 264
rect 17 260 199 263
rect 17 257 198 260
rect 17 252 196 257
rect 17 238 195 252
rect 329 249 375 277
rect 17 203 127 204
rect 17 169 35 203
rect 69 169 127 203
rect 17 127 127 169
rect 161 93 195 238
rect 17 59 35 93
rect 69 59 195 93
rect 229 209 245 243
rect 279 209 295 243
rect 229 158 295 209
rect 329 215 341 249
rect 329 198 375 215
rect 229 61 273 158
rect 409 147 443 353
rect 307 109 357 125
rect 341 75 357 109
rect 307 17 357 75
rect 391 119 443 147
rect 425 85 443 119
rect 391 51 443 85
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 397 425 431 459 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 397 85 431 119 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 213 425 247 459 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 29 153 63 187 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 235 153 269 187 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 and3_1
rlabel metal1 s 0 -48 460 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_END 3858454
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3851348
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 11.500 0.000 
<< end >>
