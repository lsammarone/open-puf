magic
tech sky130B
magscale 1 2
timestamp 1648127584
use sky130_fd_pr__hvdfm1sd2__example_55959141808719  sky130_fd_pr__hvdfm1sd2__example_55959141808719_0
timestamp 1648127584
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808719  sky130_fd_pr__hvdfm1sd2__example_55959141808719_1
timestamp 1648127584
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808719  sky130_fd_pr__hvdfm1sd2__example_55959141808719_2
timestamp 1648127584
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808782  sky130_fd_pr__hvdfm1sd__example_55959141808782_0
timestamp 1648127584
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 440 265 440 265 0 FreeSans 300 0 0 0 D
flabel comment s 284 265 284 265 0 FreeSans 300 0 0 0 S
flabel comment s 128 265 128 265 0 FreeSans 300 0 0 0 D
flabel comment s -28 265 -28 265 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 27730114
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 27728022
<< end >>
