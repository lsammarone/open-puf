magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< locali >>
rect 266 961 616 980
rect 266 855 280 961
rect 602 855 616 961
rect 266 841 616 855
rect 266 125 616 139
rect 266 19 280 125
rect 602 19 616 125
rect 266 0 616 19
<< viali >>
rect 280 855 602 961
rect 280 19 602 125
<< obsli1 >>
rect 120 817 186 883
rect 696 817 762 883
rect 120 795 160 817
rect 722 795 762 817
rect 41 759 160 795
rect 41 725 60 759
rect 94 725 160 759
rect 41 687 160 725
rect 41 653 60 687
rect 94 653 160 687
rect 41 615 160 653
rect 41 581 60 615
rect 94 581 160 615
rect 41 543 160 581
rect 41 509 60 543
rect 94 509 160 543
rect 41 471 160 509
rect 41 437 60 471
rect 94 437 160 471
rect 41 399 160 437
rect 41 365 60 399
rect 94 365 160 399
rect 41 327 160 365
rect 41 293 60 327
rect 94 293 160 327
rect 41 255 160 293
rect 41 221 60 255
rect 94 221 160 255
rect 41 185 160 221
rect 212 185 246 795
rect 318 185 352 795
rect 424 185 458 795
rect 530 185 564 795
rect 636 185 670 795
rect 722 759 841 795
rect 722 725 788 759
rect 822 725 841 759
rect 722 687 841 725
rect 722 653 788 687
rect 822 653 841 687
rect 722 615 841 653
rect 722 581 788 615
rect 822 581 841 615
rect 722 543 841 581
rect 722 509 788 543
rect 822 509 841 543
rect 722 471 841 509
rect 722 437 788 471
rect 822 437 841 471
rect 722 399 841 437
rect 722 365 788 399
rect 822 365 841 399
rect 722 327 841 365
rect 722 293 788 327
rect 822 293 841 327
rect 722 255 841 293
rect 722 221 788 255
rect 822 221 841 255
rect 722 185 841 221
rect 120 163 160 185
rect 722 163 762 185
rect 120 97 186 163
rect 696 97 762 163
<< obsli1c >>
rect 60 725 94 759
rect 60 653 94 687
rect 60 581 94 615
rect 60 509 94 543
rect 60 437 94 471
rect 60 365 94 399
rect 60 293 94 327
rect 60 221 94 255
rect 788 725 822 759
rect 788 653 822 687
rect 788 581 822 615
rect 788 509 822 543
rect 788 437 822 471
rect 788 365 822 399
rect 788 293 822 327
rect 788 221 822 255
<< metal1 >>
rect 264 961 618 980
rect 264 855 280 961
rect 602 855 618 961
rect 264 843 618 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 782 759 841 771
rect 782 725 788 759
rect 822 725 841 759
rect 782 687 841 725
rect 782 653 788 687
rect 822 653 841 687
rect 782 615 841 653
rect 782 581 788 615
rect 822 581 841 615
rect 782 543 841 581
rect 782 509 788 543
rect 822 509 841 543
rect 782 471 841 509
rect 782 437 788 471
rect 822 437 841 471
rect 782 399 841 437
rect 782 365 788 399
rect 822 365 841 399
rect 782 327 841 365
rect 782 293 788 327
rect 822 293 841 327
rect 782 255 841 293
rect 782 221 788 255
rect 822 221 841 255
rect 782 209 841 221
rect 264 125 618 137
rect 264 19 280 125
rect 602 19 618 125
rect 264 0 618 19
<< obsm1 >>
rect 203 209 255 771
rect 309 209 361 771
rect 415 209 467 771
rect 521 209 573 771
rect 627 209 679 771
<< metal2 >>
rect 14 515 868 771
rect 14 209 868 465
<< labels >>
rlabel metal2 s 14 515 868 771 6 DRAIN
port 1 nsew
rlabel viali s 280 855 602 961 6 GATE
port 2 nsew
rlabel viali s 280 19 602 125 6 GATE
port 2 nsew
rlabel locali s 266 841 616 980 6 GATE
port 2 nsew
rlabel locali s 266 0 616 139 6 GATE
port 2 nsew
rlabel metal1 s 264 843 618 980 6 GATE
port 2 nsew
rlabel metal1 s 264 0 618 137 6 GATE
port 2 nsew
rlabel metal2 s 14 209 868 465 6 SOURCE
port 3 nsew
rlabel metal1 s 41 209 100 771 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 782 209 841 771 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 14 0 868 980
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5625888
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5604998
<< end >>
