module demux2-1 (

);

endmodule
