magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< locali >>
rect 248 1369 382 1388
rect 248 1263 262 1369
rect 368 1263 382 1369
rect 248 1249 382 1263
rect 248 125 382 139
rect 248 19 262 125
rect 368 19 382 125
rect 248 0 382 19
<< viali >>
rect 262 1263 368 1369
rect 262 19 368 125
<< obsli1 >>
rect 120 1231 186 1297
rect 444 1231 510 1297
rect 120 1203 160 1231
rect 470 1203 510 1231
rect 41 1179 160 1203
rect 41 1145 60 1179
rect 94 1145 160 1179
rect 41 1107 160 1145
rect 41 1073 60 1107
rect 94 1073 160 1107
rect 41 1035 160 1073
rect 41 1001 60 1035
rect 94 1001 160 1035
rect 41 963 160 1001
rect 41 929 60 963
rect 94 929 160 963
rect 41 891 160 929
rect 41 857 60 891
rect 94 857 160 891
rect 41 819 160 857
rect 41 785 60 819
rect 94 785 160 819
rect 41 747 160 785
rect 41 713 60 747
rect 94 713 160 747
rect 41 675 160 713
rect 41 641 60 675
rect 94 641 160 675
rect 41 603 160 641
rect 41 569 60 603
rect 94 569 160 603
rect 41 531 160 569
rect 41 497 60 531
rect 94 497 160 531
rect 41 459 160 497
rect 41 425 60 459
rect 94 425 160 459
rect 41 387 160 425
rect 41 353 60 387
rect 94 353 160 387
rect 41 315 160 353
rect 41 281 60 315
rect 94 281 160 315
rect 41 243 160 281
rect 41 209 60 243
rect 94 209 160 243
rect 41 185 160 209
rect 212 185 246 1203
rect 298 185 332 1203
rect 384 185 418 1203
rect 470 1179 589 1203
rect 470 1145 536 1179
rect 570 1145 589 1179
rect 470 1107 589 1145
rect 470 1073 536 1107
rect 570 1073 589 1107
rect 470 1035 589 1073
rect 470 1001 536 1035
rect 570 1001 589 1035
rect 470 963 589 1001
rect 470 929 536 963
rect 570 929 589 963
rect 470 891 589 929
rect 470 857 536 891
rect 570 857 589 891
rect 470 819 589 857
rect 470 785 536 819
rect 570 785 589 819
rect 470 747 589 785
rect 470 713 536 747
rect 570 713 589 747
rect 470 675 589 713
rect 470 641 536 675
rect 570 641 589 675
rect 470 603 589 641
rect 470 569 536 603
rect 570 569 589 603
rect 470 531 589 569
rect 470 497 536 531
rect 570 497 589 531
rect 470 459 589 497
rect 470 425 536 459
rect 570 425 589 459
rect 470 387 589 425
rect 470 353 536 387
rect 570 353 589 387
rect 470 315 589 353
rect 470 281 536 315
rect 570 281 589 315
rect 470 243 589 281
rect 470 209 536 243
rect 570 209 589 243
rect 470 185 589 209
rect 120 157 160 185
rect 470 157 510 185
rect 120 91 186 157
rect 444 91 510 157
<< obsli1c >>
rect 60 1145 94 1179
rect 60 1073 94 1107
rect 60 1001 94 1035
rect 60 929 94 963
rect 60 857 94 891
rect 60 785 94 819
rect 60 713 94 747
rect 60 641 94 675
rect 60 569 94 603
rect 60 497 94 531
rect 60 425 94 459
rect 60 353 94 387
rect 60 281 94 315
rect 60 209 94 243
rect 536 1145 570 1179
rect 536 1073 570 1107
rect 536 1001 570 1035
rect 536 929 570 963
rect 536 857 570 891
rect 536 785 570 819
rect 536 713 570 747
rect 536 641 570 675
rect 536 569 570 603
rect 536 497 570 531
rect 536 425 570 459
rect 536 353 570 387
rect 536 281 570 315
rect 536 209 570 243
<< metal1 >>
rect 250 1369 380 1388
rect 250 1263 262 1369
rect 368 1263 380 1369
rect 250 1251 380 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 530 1179 589 1191
rect 530 1145 536 1179
rect 570 1145 589 1179
rect 530 1107 589 1145
rect 530 1073 536 1107
rect 570 1073 589 1107
rect 530 1035 589 1073
rect 530 1001 536 1035
rect 570 1001 589 1035
rect 530 963 589 1001
rect 530 929 536 963
rect 570 929 589 963
rect 530 891 589 929
rect 530 857 536 891
rect 570 857 589 891
rect 530 819 589 857
rect 530 785 536 819
rect 570 785 589 819
rect 530 747 589 785
rect 530 713 536 747
rect 570 713 589 747
rect 530 675 589 713
rect 530 641 536 675
rect 570 641 589 675
rect 530 603 589 641
rect 530 569 536 603
rect 570 569 589 603
rect 530 531 589 569
rect 530 497 536 531
rect 570 497 589 531
rect 530 459 589 497
rect 530 425 536 459
rect 570 425 589 459
rect 530 387 589 425
rect 530 353 536 387
rect 570 353 589 387
rect 530 315 589 353
rect 530 281 536 315
rect 570 281 589 315
rect 530 243 589 281
rect 530 209 536 243
rect 570 209 589 243
rect 530 197 589 209
rect 250 125 380 137
rect 250 19 262 125
rect 368 19 380 125
rect 250 0 380 19
<< obsm1 >>
rect 203 197 255 1191
rect 289 197 341 1191
rect 375 197 427 1191
<< metal2 >>
rect 14 719 616 1191
rect 14 197 616 669
<< labels >>
rlabel metal1 s 530 197 589 1191 6 BULK
port 1 nsew
rlabel metal1 s 41 197 100 1191 6 BULK
port 1 nsew
rlabel metal2 s 14 719 616 1191 6 DRAIN
port 2 nsew
rlabel viali s 262 1263 368 1369 6 GATE
port 3 nsew
rlabel viali s 262 19 368 125 6 GATE
port 3 nsew
rlabel locali s 248 1249 382 1388 6 GATE
port 3 nsew
rlabel locali s 248 0 382 139 6 GATE
port 3 nsew
rlabel metal1 s 250 1251 380 1388 6 GATE
port 3 nsew
rlabel metal1 s 250 0 380 137 6 GATE
port 3 nsew
rlabel metal2 s 14 197 616 669 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 630 1388
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9851430
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9831346
<< end >>
