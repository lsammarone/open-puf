magic
tech sky130A
magscale 1 2
timestamp 1648127584
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_0
timestamp 1648127584
transform 1 0 581 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_1
timestamp 1648127584
transform 1 0 1501 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_2
timestamp 1648127584
transform 1 0 2421 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_3
timestamp 1648127584
transform 1 0 3341 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_4
timestamp 1648127584
transform 1 0 4261 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_5
timestamp 1648127584
transform 1 0 5181 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_6
timestamp 1648127584
transform 1 0 6101 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_7
timestamp 1648127584
transform 1 0 7021 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_8
timestamp 1648127584
transform 1 0 7941 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808676  sky130_fd_pr__hvdftpl1s2__example_55959141808676_9
timestamp 1648127584
transform 1 0 8861 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s__example_55959141808675  sky130_fd_pr__hvdftpl1s__example_55959141808675_0
timestamp 1648127584
transform -1 0 -79 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s__example_55959141808675  sky130_fd_pr__hvdftpl1s__example_55959141808675_1
timestamp 1648127584
transform 1 0 9781 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 9843 987 9843 987 0 FreeSans 300 0 0 0 S
flabel comment s 9451 1000 9451 1000 0 FreeSans 300 0 0 0 D
flabel comment s 8991 981 8991 981 0 FreeSans 300 0 0 0 S
flabel comment s 8531 1000 8531 1000 0 FreeSans 300 0 0 0 D
flabel comment s 8071 981 8071 981 0 FreeSans 300 0 0 0 S
flabel comment s 7611 1000 7611 1000 0 FreeSans 300 0 0 0 D
flabel comment s 7151 981 7151 981 0 FreeSans 300 0 0 0 S
flabel comment s 6691 1000 6691 1000 0 FreeSans 300 0 0 0 D
flabel comment s 6231 981 6231 981 0 FreeSans 300 0 0 0 S
flabel comment s 5771 1000 5771 1000 0 FreeSans 300 0 0 0 D
flabel comment s 5311 981 5311 981 0 FreeSans 300 0 0 0 S
flabel comment s 4851 1000 4851 1000 0 FreeSans 300 0 0 0 D
flabel comment s 4391 981 4391 981 0 FreeSans 300 0 0 0 S
flabel comment s 3931 1000 3931 1000 0 FreeSans 300 0 0 0 D
flabel comment s 3471 981 3471 981 0 FreeSans 300 0 0 0 S
flabel comment s 3011 1000 3011 1000 0 FreeSans 300 0 0 0 D
flabel comment s 2551 981 2551 981 0 FreeSans 300 0 0 0 S
flabel comment s 2091 1000 2091 1000 0 FreeSans 300 0 0 0 D
flabel comment s 1631 981 1631 981 0 FreeSans 300 0 0 0 S
flabel comment s 1171 1000 1171 1000 0 FreeSans 300 0 0 0 D
flabel comment s 711 981 711 981 0 FreeSans 300 0 0 0 S
flabel comment s 251 1000 251 1000 0 FreeSans 300 0 0 0 D
flabel comment s -141 987 -141 987 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 11221224
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 11209504
<< end >>
