magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 314 582
<< pwell >>
rect 1 21 275 177
rect 213 -17 247 21
<< locali >>
rect 17 312 71 493
rect 17 152 51 312
rect 189 197 255 271
rect 17 51 69 152
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 105 459 171 493
rect 105 425 122 459
rect 156 425 171 459
rect 105 375 171 425
rect 207 341 241 493
rect 108 307 241 341
rect 108 278 142 307
rect 85 212 142 278
rect 108 161 142 212
rect 108 127 241 161
rect 105 17 171 93
rect 207 51 241 127
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 122 425 156 459
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
<< metal1 >>
rect 0 561 276 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 276 561
rect 0 496 276 527
rect 14 459 262 468
rect 14 428 122 459
rect 110 425 122 428
rect 156 428 262 459
rect 156 425 168 428
rect 110 416 168 425
rect 0 17 276 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 276 17
rect 0 -48 276 -17
<< labels >>
rlabel locali s 189 197 255 271 6 A
port 1 nsew signal input
rlabel metal1 s 110 416 168 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 14 428 262 468 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 -48 276 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 213 -17 247 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 275 177 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 314 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 276 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 17 51 69 152 6 X
port 7 nsew signal output
rlabel locali s 17 152 51 312 6 X
port 7 nsew signal output
rlabel locali s 17 312 71 493 6 X
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 276 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2180928
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2176844
<< end >>
