magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 1 21 459 203
rect 29 -17 63 21
<< locali >>
rect 18 333 85 490
rect 18 299 135 333
rect 206 323 257 490
rect 17 149 67 265
rect 101 165 135 299
rect 169 283 257 323
rect 169 199 215 283
rect 291 249 339 490
rect 249 215 339 249
rect 101 131 341 165
rect 391 131 443 333
rect 101 129 172 131
rect 119 77 172 129
rect 307 77 341 131
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 391 367 443 527
rect 17 17 69 115
rect 207 17 273 97
rect 375 17 441 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 391 131 443 333 6 A
port 1 nsew signal input
rlabel locali s 249 215 339 249 6 B
port 2 nsew signal input
rlabel locali s 291 249 339 490 6 B
port 2 nsew signal input
rlabel locali s 169 199 215 283 6 C
port 3 nsew signal input
rlabel locali s 169 283 257 323 6 C
port 3 nsew signal input
rlabel locali s 206 323 257 490 6 C
port 3 nsew signal input
rlabel locali s 17 149 67 265 6 D
port 4 nsew signal input
rlabel metal1 s 0 -48 460 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 459 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 307 77 341 131 6 Y
port 9 nsew signal output
rlabel locali s 119 77 172 129 6 Y
port 9 nsew signal output
rlabel locali s 101 129 172 131 6 Y
port 9 nsew signal output
rlabel locali s 101 131 341 165 6 Y
port 9 nsew signal output
rlabel locali s 101 165 135 299 6 Y
port 9 nsew signal output
rlabel locali s 18 299 135 333 6 Y
port 9 nsew signal output
rlabel locali s 18 333 85 490 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 460 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1151400
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1146680
<< end >>
