/farmshare/home/classes/ee/372/PDKs/share/pdk/sky130A/libs.tech/ngspice/sonos_see_p/begin_of_life/typical.spice