magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< obsli1 >>
rect 26 669 770 770
rect 26 127 127 669
rect 189 535 607 607
rect 189 261 261 535
rect 319 319 477 477
rect 535 261 607 535
rect 189 189 607 261
rect 669 127 770 669
rect 26 26 770 127
<< obsm1 >>
rect 315 315 481 481
<< properties >>
string FIXED_BBOX 26 26 770 795
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3986574
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 3979106
<< end >>
