magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -1 766 3131 892
rect 3149 766 6281 892
rect 6299 766 9431 1334
rect 9449 766 12581 1334
rect 12599 766 15731 1334
rect 15749 766 18881 1334
rect 18899 766 22031 1334
rect 22274 766 24406 2180
rect -1 554 24406 766
rect 6299 528 9431 554
rect 9449 528 12581 554
rect 12599 528 15731 554
rect 15749 528 18881 554
rect 18899 528 22031 554
<< mvpmos >>
rect 22340 1961 24340 2061
rect 22340 1805 24340 1905
rect 22340 1649 24340 1749
rect 22340 1493 24340 1593
rect 22340 1337 24340 1437
rect 6365 1115 9365 1215
rect 9515 1115 12515 1215
rect 12665 1115 15665 1215
rect 15815 1115 18815 1215
rect 18965 1115 21965 1215
rect 6365 959 9365 1059
rect 9515 959 12515 1059
rect 65 673 3065 773
rect 6365 803 9365 903
rect 12665 959 15665 1059
rect 9515 803 12515 903
rect 15815 959 18815 1059
rect 12665 803 15665 903
rect 18965 959 21965 1059
rect 15815 803 18815 903
rect 18965 803 21965 903
rect 3215 673 6215 773
rect 6365 647 9365 747
rect 9515 647 12515 747
rect 12665 647 15665 747
rect 15815 647 18815 747
rect 18965 647 21965 747
rect 22340 1181 24340 1281
rect 22340 1025 24340 1125
rect 22340 869 24340 969
rect 22340 713 24340 813
<< mvpdiff >>
rect 22340 2106 24340 2114
rect 22340 2072 22390 2106
rect 22424 2072 22458 2106
rect 22492 2072 22526 2106
rect 22560 2072 22594 2106
rect 22628 2072 22662 2106
rect 22696 2072 22730 2106
rect 22764 2072 22798 2106
rect 22832 2072 22866 2106
rect 22900 2072 22934 2106
rect 22968 2072 23002 2106
rect 23036 2072 23070 2106
rect 23104 2072 23138 2106
rect 23172 2072 23206 2106
rect 23240 2072 23274 2106
rect 23308 2072 23342 2106
rect 23376 2072 23410 2106
rect 23444 2072 23478 2106
rect 23512 2072 23546 2106
rect 23580 2072 23614 2106
rect 23648 2072 23682 2106
rect 23716 2072 23750 2106
rect 23784 2072 23818 2106
rect 23852 2072 23886 2106
rect 23920 2072 23954 2106
rect 23988 2072 24022 2106
rect 24056 2072 24090 2106
rect 24124 2072 24158 2106
rect 24192 2072 24226 2106
rect 24260 2072 24294 2106
rect 24328 2072 24340 2106
rect 22340 2061 24340 2072
rect 22340 1950 24340 1961
rect 22340 1916 22390 1950
rect 22424 1916 22458 1950
rect 22492 1916 22526 1950
rect 22560 1916 22594 1950
rect 22628 1916 22662 1950
rect 22696 1916 22730 1950
rect 22764 1916 22798 1950
rect 22832 1916 22866 1950
rect 22900 1916 22934 1950
rect 22968 1916 23002 1950
rect 23036 1916 23070 1950
rect 23104 1916 23138 1950
rect 23172 1916 23206 1950
rect 23240 1916 23274 1950
rect 23308 1916 23342 1950
rect 23376 1916 23410 1950
rect 23444 1916 23478 1950
rect 23512 1916 23546 1950
rect 23580 1916 23614 1950
rect 23648 1916 23682 1950
rect 23716 1916 23750 1950
rect 23784 1916 23818 1950
rect 23852 1916 23886 1950
rect 23920 1916 23954 1950
rect 23988 1916 24022 1950
rect 24056 1916 24090 1950
rect 24124 1916 24158 1950
rect 24192 1916 24226 1950
rect 24260 1916 24294 1950
rect 24328 1916 24340 1950
rect 22340 1905 24340 1916
rect 22340 1794 24340 1805
rect 22340 1760 22390 1794
rect 22424 1760 22458 1794
rect 22492 1760 22526 1794
rect 22560 1760 22594 1794
rect 22628 1760 22662 1794
rect 22696 1760 22730 1794
rect 22764 1760 22798 1794
rect 22832 1760 22866 1794
rect 22900 1760 22934 1794
rect 22968 1760 23002 1794
rect 23036 1760 23070 1794
rect 23104 1760 23138 1794
rect 23172 1760 23206 1794
rect 23240 1760 23274 1794
rect 23308 1760 23342 1794
rect 23376 1760 23410 1794
rect 23444 1760 23478 1794
rect 23512 1760 23546 1794
rect 23580 1760 23614 1794
rect 23648 1760 23682 1794
rect 23716 1760 23750 1794
rect 23784 1760 23818 1794
rect 23852 1760 23886 1794
rect 23920 1760 23954 1794
rect 23988 1760 24022 1794
rect 24056 1760 24090 1794
rect 24124 1760 24158 1794
rect 24192 1760 24226 1794
rect 24260 1760 24294 1794
rect 24328 1760 24340 1794
rect 22340 1749 24340 1760
rect 22340 1638 24340 1649
rect 22340 1604 22390 1638
rect 22424 1604 22458 1638
rect 22492 1604 22526 1638
rect 22560 1604 22594 1638
rect 22628 1604 22662 1638
rect 22696 1604 22730 1638
rect 22764 1604 22798 1638
rect 22832 1604 22866 1638
rect 22900 1604 22934 1638
rect 22968 1604 23002 1638
rect 23036 1604 23070 1638
rect 23104 1604 23138 1638
rect 23172 1604 23206 1638
rect 23240 1604 23274 1638
rect 23308 1604 23342 1638
rect 23376 1604 23410 1638
rect 23444 1604 23478 1638
rect 23512 1604 23546 1638
rect 23580 1604 23614 1638
rect 23648 1604 23682 1638
rect 23716 1604 23750 1638
rect 23784 1604 23818 1638
rect 23852 1604 23886 1638
rect 23920 1604 23954 1638
rect 23988 1604 24022 1638
rect 24056 1604 24090 1638
rect 24124 1604 24158 1638
rect 24192 1604 24226 1638
rect 24260 1604 24294 1638
rect 24328 1604 24340 1638
rect 22340 1593 24340 1604
rect 22340 1482 24340 1493
rect 22340 1448 22390 1482
rect 22424 1448 22458 1482
rect 22492 1448 22526 1482
rect 22560 1448 22594 1482
rect 22628 1448 22662 1482
rect 22696 1448 22730 1482
rect 22764 1448 22798 1482
rect 22832 1448 22866 1482
rect 22900 1448 22934 1482
rect 22968 1448 23002 1482
rect 23036 1448 23070 1482
rect 23104 1448 23138 1482
rect 23172 1448 23206 1482
rect 23240 1448 23274 1482
rect 23308 1448 23342 1482
rect 23376 1448 23410 1482
rect 23444 1448 23478 1482
rect 23512 1448 23546 1482
rect 23580 1448 23614 1482
rect 23648 1448 23682 1482
rect 23716 1448 23750 1482
rect 23784 1448 23818 1482
rect 23852 1448 23886 1482
rect 23920 1448 23954 1482
rect 23988 1448 24022 1482
rect 24056 1448 24090 1482
rect 24124 1448 24158 1482
rect 24192 1448 24226 1482
rect 24260 1448 24294 1482
rect 24328 1448 24340 1482
rect 22340 1437 24340 1448
rect 22340 1326 24340 1337
rect 22340 1292 22390 1326
rect 22424 1292 22458 1326
rect 22492 1292 22526 1326
rect 22560 1292 22594 1326
rect 22628 1292 22662 1326
rect 22696 1292 22730 1326
rect 22764 1292 22798 1326
rect 22832 1292 22866 1326
rect 22900 1292 22934 1326
rect 22968 1292 23002 1326
rect 23036 1292 23070 1326
rect 23104 1292 23138 1326
rect 23172 1292 23206 1326
rect 23240 1292 23274 1326
rect 23308 1292 23342 1326
rect 23376 1292 23410 1326
rect 23444 1292 23478 1326
rect 23512 1292 23546 1326
rect 23580 1292 23614 1326
rect 23648 1292 23682 1326
rect 23716 1292 23750 1326
rect 23784 1292 23818 1326
rect 23852 1292 23886 1326
rect 23920 1292 23954 1326
rect 23988 1292 24022 1326
rect 24056 1292 24090 1326
rect 24124 1292 24158 1326
rect 24192 1292 24226 1326
rect 24260 1292 24294 1326
rect 24328 1292 24340 1326
rect 22340 1281 24340 1292
rect 6365 1260 9365 1268
rect 6365 1226 6395 1260
rect 6429 1226 6463 1260
rect 6497 1226 6531 1260
rect 6565 1226 6599 1260
rect 6633 1226 6667 1260
rect 6701 1226 6735 1260
rect 6769 1226 6803 1260
rect 6837 1226 6871 1260
rect 6905 1226 6939 1260
rect 6973 1226 7007 1260
rect 7041 1226 7075 1260
rect 7109 1226 7143 1260
rect 7177 1226 7211 1260
rect 7245 1226 7279 1260
rect 7313 1226 7347 1260
rect 7381 1226 7415 1260
rect 7449 1226 7483 1260
rect 7517 1226 7551 1260
rect 7585 1226 7619 1260
rect 7653 1226 7687 1260
rect 7721 1226 7755 1260
rect 7789 1226 7823 1260
rect 7857 1226 7891 1260
rect 7925 1226 7959 1260
rect 7993 1226 8027 1260
rect 8061 1226 8095 1260
rect 8129 1226 8163 1260
rect 8197 1226 8231 1260
rect 8265 1226 8299 1260
rect 8333 1226 8367 1260
rect 8401 1226 8435 1260
rect 8469 1226 8503 1260
rect 8537 1226 8571 1260
rect 8605 1226 8639 1260
rect 8673 1226 8707 1260
rect 8741 1226 8775 1260
rect 8809 1226 8843 1260
rect 8877 1226 8911 1260
rect 8945 1226 8979 1260
rect 9013 1226 9047 1260
rect 9081 1226 9115 1260
rect 9149 1226 9183 1260
rect 9217 1226 9251 1260
rect 9285 1226 9319 1260
rect 9353 1226 9365 1260
rect 6365 1215 9365 1226
rect 9515 1260 12515 1268
rect 9515 1226 9545 1260
rect 9579 1226 9613 1260
rect 9647 1226 9681 1260
rect 9715 1226 9749 1260
rect 9783 1226 9817 1260
rect 9851 1226 9885 1260
rect 9919 1226 9953 1260
rect 9987 1226 10021 1260
rect 10055 1226 10089 1260
rect 10123 1226 10157 1260
rect 10191 1226 10225 1260
rect 10259 1226 10293 1260
rect 10327 1226 10361 1260
rect 10395 1226 10429 1260
rect 10463 1226 10497 1260
rect 10531 1226 10565 1260
rect 10599 1226 10633 1260
rect 10667 1226 10701 1260
rect 10735 1226 10769 1260
rect 10803 1226 10837 1260
rect 10871 1226 10905 1260
rect 10939 1226 10973 1260
rect 11007 1226 11041 1260
rect 11075 1226 11109 1260
rect 11143 1226 11177 1260
rect 11211 1226 11245 1260
rect 11279 1226 11313 1260
rect 11347 1226 11381 1260
rect 11415 1226 11449 1260
rect 11483 1226 11517 1260
rect 11551 1226 11585 1260
rect 11619 1226 11653 1260
rect 11687 1226 11721 1260
rect 11755 1226 11789 1260
rect 11823 1226 11857 1260
rect 11891 1226 11925 1260
rect 11959 1226 11993 1260
rect 12027 1226 12061 1260
rect 12095 1226 12129 1260
rect 12163 1226 12197 1260
rect 12231 1226 12265 1260
rect 12299 1226 12333 1260
rect 12367 1226 12401 1260
rect 12435 1226 12469 1260
rect 12503 1226 12515 1260
rect 9515 1215 12515 1226
rect 12665 1260 15665 1268
rect 12665 1226 12695 1260
rect 12729 1226 12763 1260
rect 12797 1226 12831 1260
rect 12865 1226 12899 1260
rect 12933 1226 12967 1260
rect 13001 1226 13035 1260
rect 13069 1226 13103 1260
rect 13137 1226 13171 1260
rect 13205 1226 13239 1260
rect 13273 1226 13307 1260
rect 13341 1226 13375 1260
rect 13409 1226 13443 1260
rect 13477 1226 13511 1260
rect 13545 1226 13579 1260
rect 13613 1226 13647 1260
rect 13681 1226 13715 1260
rect 13749 1226 13783 1260
rect 13817 1226 13851 1260
rect 13885 1226 13919 1260
rect 13953 1226 13987 1260
rect 14021 1226 14055 1260
rect 14089 1226 14123 1260
rect 14157 1226 14191 1260
rect 14225 1226 14259 1260
rect 14293 1226 14327 1260
rect 14361 1226 14395 1260
rect 14429 1226 14463 1260
rect 14497 1226 14531 1260
rect 14565 1226 14599 1260
rect 14633 1226 14667 1260
rect 14701 1226 14735 1260
rect 14769 1226 14803 1260
rect 14837 1226 14871 1260
rect 14905 1226 14939 1260
rect 14973 1226 15007 1260
rect 15041 1226 15075 1260
rect 15109 1226 15143 1260
rect 15177 1226 15211 1260
rect 15245 1226 15279 1260
rect 15313 1226 15347 1260
rect 15381 1226 15415 1260
rect 15449 1226 15483 1260
rect 15517 1226 15551 1260
rect 15585 1226 15619 1260
rect 15653 1226 15665 1260
rect 12665 1215 15665 1226
rect 15815 1260 18815 1268
rect 15815 1226 15845 1260
rect 15879 1226 15913 1260
rect 15947 1226 15981 1260
rect 16015 1226 16049 1260
rect 16083 1226 16117 1260
rect 16151 1226 16185 1260
rect 16219 1226 16253 1260
rect 16287 1226 16321 1260
rect 16355 1226 16389 1260
rect 16423 1226 16457 1260
rect 16491 1226 16525 1260
rect 16559 1226 16593 1260
rect 16627 1226 16661 1260
rect 16695 1226 16729 1260
rect 16763 1226 16797 1260
rect 16831 1226 16865 1260
rect 16899 1226 16933 1260
rect 16967 1226 17001 1260
rect 17035 1226 17069 1260
rect 17103 1226 17137 1260
rect 17171 1226 17205 1260
rect 17239 1226 17273 1260
rect 17307 1226 17341 1260
rect 17375 1226 17409 1260
rect 17443 1226 17477 1260
rect 17511 1226 17545 1260
rect 17579 1226 17613 1260
rect 17647 1226 17681 1260
rect 17715 1226 17749 1260
rect 17783 1226 17817 1260
rect 17851 1226 17885 1260
rect 17919 1226 17953 1260
rect 17987 1226 18021 1260
rect 18055 1226 18089 1260
rect 18123 1226 18157 1260
rect 18191 1226 18225 1260
rect 18259 1226 18293 1260
rect 18327 1226 18361 1260
rect 18395 1226 18429 1260
rect 18463 1226 18497 1260
rect 18531 1226 18565 1260
rect 18599 1226 18633 1260
rect 18667 1226 18701 1260
rect 18735 1226 18769 1260
rect 18803 1226 18815 1260
rect 15815 1215 18815 1226
rect 18965 1260 21965 1268
rect 18965 1226 18995 1260
rect 19029 1226 19063 1260
rect 19097 1226 19131 1260
rect 19165 1226 19199 1260
rect 19233 1226 19267 1260
rect 19301 1226 19335 1260
rect 19369 1226 19403 1260
rect 19437 1226 19471 1260
rect 19505 1226 19539 1260
rect 19573 1226 19607 1260
rect 19641 1226 19675 1260
rect 19709 1226 19743 1260
rect 19777 1226 19811 1260
rect 19845 1226 19879 1260
rect 19913 1226 19947 1260
rect 19981 1226 20015 1260
rect 20049 1226 20083 1260
rect 20117 1226 20151 1260
rect 20185 1226 20219 1260
rect 20253 1226 20287 1260
rect 20321 1226 20355 1260
rect 20389 1226 20423 1260
rect 20457 1226 20491 1260
rect 20525 1226 20559 1260
rect 20593 1226 20627 1260
rect 20661 1226 20695 1260
rect 20729 1226 20763 1260
rect 20797 1226 20831 1260
rect 20865 1226 20899 1260
rect 20933 1226 20967 1260
rect 21001 1226 21035 1260
rect 21069 1226 21103 1260
rect 21137 1226 21171 1260
rect 21205 1226 21239 1260
rect 21273 1226 21307 1260
rect 21341 1226 21375 1260
rect 21409 1226 21443 1260
rect 21477 1226 21511 1260
rect 21545 1226 21579 1260
rect 21613 1226 21647 1260
rect 21681 1226 21715 1260
rect 21749 1226 21783 1260
rect 21817 1226 21851 1260
rect 21885 1226 21919 1260
rect 21953 1226 21965 1260
rect 18965 1215 21965 1226
rect 6365 1104 9365 1115
rect 6365 1070 6395 1104
rect 6429 1070 6463 1104
rect 6497 1070 6531 1104
rect 6565 1070 6599 1104
rect 6633 1070 6667 1104
rect 6701 1070 6735 1104
rect 6769 1070 6803 1104
rect 6837 1070 6871 1104
rect 6905 1070 6939 1104
rect 6973 1070 7007 1104
rect 7041 1070 7075 1104
rect 7109 1070 7143 1104
rect 7177 1070 7211 1104
rect 7245 1070 7279 1104
rect 7313 1070 7347 1104
rect 7381 1070 7415 1104
rect 7449 1070 7483 1104
rect 7517 1070 7551 1104
rect 7585 1070 7619 1104
rect 7653 1070 7687 1104
rect 7721 1070 7755 1104
rect 7789 1070 7823 1104
rect 7857 1070 7891 1104
rect 7925 1070 7959 1104
rect 7993 1070 8027 1104
rect 8061 1070 8095 1104
rect 8129 1070 8163 1104
rect 8197 1070 8231 1104
rect 8265 1070 8299 1104
rect 8333 1070 8367 1104
rect 8401 1070 8435 1104
rect 8469 1070 8503 1104
rect 8537 1070 8571 1104
rect 8605 1070 8639 1104
rect 8673 1070 8707 1104
rect 8741 1070 8775 1104
rect 8809 1070 8843 1104
rect 8877 1070 8911 1104
rect 8945 1070 8979 1104
rect 9013 1070 9047 1104
rect 9081 1070 9115 1104
rect 9149 1070 9183 1104
rect 9217 1070 9251 1104
rect 9285 1070 9319 1104
rect 9353 1070 9365 1104
rect 6365 1059 9365 1070
rect 9515 1104 12515 1115
rect 9515 1070 9545 1104
rect 9579 1070 9613 1104
rect 9647 1070 9681 1104
rect 9715 1070 9749 1104
rect 9783 1070 9817 1104
rect 9851 1070 9885 1104
rect 9919 1070 9953 1104
rect 9987 1070 10021 1104
rect 10055 1070 10089 1104
rect 10123 1070 10157 1104
rect 10191 1070 10225 1104
rect 10259 1070 10293 1104
rect 10327 1070 10361 1104
rect 10395 1070 10429 1104
rect 10463 1070 10497 1104
rect 10531 1070 10565 1104
rect 10599 1070 10633 1104
rect 10667 1070 10701 1104
rect 10735 1070 10769 1104
rect 10803 1070 10837 1104
rect 10871 1070 10905 1104
rect 10939 1070 10973 1104
rect 11007 1070 11041 1104
rect 11075 1070 11109 1104
rect 11143 1070 11177 1104
rect 11211 1070 11245 1104
rect 11279 1070 11313 1104
rect 11347 1070 11381 1104
rect 11415 1070 11449 1104
rect 11483 1070 11517 1104
rect 11551 1070 11585 1104
rect 11619 1070 11653 1104
rect 11687 1070 11721 1104
rect 11755 1070 11789 1104
rect 11823 1070 11857 1104
rect 11891 1070 11925 1104
rect 11959 1070 11993 1104
rect 12027 1070 12061 1104
rect 12095 1070 12129 1104
rect 12163 1070 12197 1104
rect 12231 1070 12265 1104
rect 12299 1070 12333 1104
rect 12367 1070 12401 1104
rect 12435 1070 12469 1104
rect 12503 1070 12515 1104
rect 9515 1059 12515 1070
rect 12665 1104 15665 1115
rect 12665 1070 12695 1104
rect 12729 1070 12763 1104
rect 12797 1070 12831 1104
rect 12865 1070 12899 1104
rect 12933 1070 12967 1104
rect 13001 1070 13035 1104
rect 13069 1070 13103 1104
rect 13137 1070 13171 1104
rect 13205 1070 13239 1104
rect 13273 1070 13307 1104
rect 13341 1070 13375 1104
rect 13409 1070 13443 1104
rect 13477 1070 13511 1104
rect 13545 1070 13579 1104
rect 13613 1070 13647 1104
rect 13681 1070 13715 1104
rect 13749 1070 13783 1104
rect 13817 1070 13851 1104
rect 13885 1070 13919 1104
rect 13953 1070 13987 1104
rect 14021 1070 14055 1104
rect 14089 1070 14123 1104
rect 14157 1070 14191 1104
rect 14225 1070 14259 1104
rect 14293 1070 14327 1104
rect 14361 1070 14395 1104
rect 14429 1070 14463 1104
rect 14497 1070 14531 1104
rect 14565 1070 14599 1104
rect 14633 1070 14667 1104
rect 14701 1070 14735 1104
rect 14769 1070 14803 1104
rect 14837 1070 14871 1104
rect 14905 1070 14939 1104
rect 14973 1070 15007 1104
rect 15041 1070 15075 1104
rect 15109 1070 15143 1104
rect 15177 1070 15211 1104
rect 15245 1070 15279 1104
rect 15313 1070 15347 1104
rect 15381 1070 15415 1104
rect 15449 1070 15483 1104
rect 15517 1070 15551 1104
rect 15585 1070 15619 1104
rect 15653 1070 15665 1104
rect 12665 1059 15665 1070
rect 15815 1104 18815 1115
rect 15815 1070 15845 1104
rect 15879 1070 15913 1104
rect 15947 1070 15981 1104
rect 16015 1070 16049 1104
rect 16083 1070 16117 1104
rect 16151 1070 16185 1104
rect 16219 1070 16253 1104
rect 16287 1070 16321 1104
rect 16355 1070 16389 1104
rect 16423 1070 16457 1104
rect 16491 1070 16525 1104
rect 16559 1070 16593 1104
rect 16627 1070 16661 1104
rect 16695 1070 16729 1104
rect 16763 1070 16797 1104
rect 16831 1070 16865 1104
rect 16899 1070 16933 1104
rect 16967 1070 17001 1104
rect 17035 1070 17069 1104
rect 17103 1070 17137 1104
rect 17171 1070 17205 1104
rect 17239 1070 17273 1104
rect 17307 1070 17341 1104
rect 17375 1070 17409 1104
rect 17443 1070 17477 1104
rect 17511 1070 17545 1104
rect 17579 1070 17613 1104
rect 17647 1070 17681 1104
rect 17715 1070 17749 1104
rect 17783 1070 17817 1104
rect 17851 1070 17885 1104
rect 17919 1070 17953 1104
rect 17987 1070 18021 1104
rect 18055 1070 18089 1104
rect 18123 1070 18157 1104
rect 18191 1070 18225 1104
rect 18259 1070 18293 1104
rect 18327 1070 18361 1104
rect 18395 1070 18429 1104
rect 18463 1070 18497 1104
rect 18531 1070 18565 1104
rect 18599 1070 18633 1104
rect 18667 1070 18701 1104
rect 18735 1070 18769 1104
rect 18803 1070 18815 1104
rect 15815 1059 18815 1070
rect 18965 1104 21965 1115
rect 18965 1070 18995 1104
rect 19029 1070 19063 1104
rect 19097 1070 19131 1104
rect 19165 1070 19199 1104
rect 19233 1070 19267 1104
rect 19301 1070 19335 1104
rect 19369 1070 19403 1104
rect 19437 1070 19471 1104
rect 19505 1070 19539 1104
rect 19573 1070 19607 1104
rect 19641 1070 19675 1104
rect 19709 1070 19743 1104
rect 19777 1070 19811 1104
rect 19845 1070 19879 1104
rect 19913 1070 19947 1104
rect 19981 1070 20015 1104
rect 20049 1070 20083 1104
rect 20117 1070 20151 1104
rect 20185 1070 20219 1104
rect 20253 1070 20287 1104
rect 20321 1070 20355 1104
rect 20389 1070 20423 1104
rect 20457 1070 20491 1104
rect 20525 1070 20559 1104
rect 20593 1070 20627 1104
rect 20661 1070 20695 1104
rect 20729 1070 20763 1104
rect 20797 1070 20831 1104
rect 20865 1070 20899 1104
rect 20933 1070 20967 1104
rect 21001 1070 21035 1104
rect 21069 1070 21103 1104
rect 21137 1070 21171 1104
rect 21205 1070 21239 1104
rect 21273 1070 21307 1104
rect 21341 1070 21375 1104
rect 21409 1070 21443 1104
rect 21477 1070 21511 1104
rect 21545 1070 21579 1104
rect 21613 1070 21647 1104
rect 21681 1070 21715 1104
rect 21749 1070 21783 1104
rect 21817 1070 21851 1104
rect 21885 1070 21919 1104
rect 21953 1070 21965 1104
rect 18965 1059 21965 1070
rect 6365 948 9365 959
rect 6365 914 6395 948
rect 6429 914 6463 948
rect 6497 914 6531 948
rect 6565 914 6599 948
rect 6633 914 6667 948
rect 6701 914 6735 948
rect 6769 914 6803 948
rect 6837 914 6871 948
rect 6905 914 6939 948
rect 6973 914 7007 948
rect 7041 914 7075 948
rect 7109 914 7143 948
rect 7177 914 7211 948
rect 7245 914 7279 948
rect 7313 914 7347 948
rect 7381 914 7415 948
rect 7449 914 7483 948
rect 7517 914 7551 948
rect 7585 914 7619 948
rect 7653 914 7687 948
rect 7721 914 7755 948
rect 7789 914 7823 948
rect 7857 914 7891 948
rect 7925 914 7959 948
rect 7993 914 8027 948
rect 8061 914 8095 948
rect 8129 914 8163 948
rect 8197 914 8231 948
rect 8265 914 8299 948
rect 8333 914 8367 948
rect 8401 914 8435 948
rect 8469 914 8503 948
rect 8537 914 8571 948
rect 8605 914 8639 948
rect 8673 914 8707 948
rect 8741 914 8775 948
rect 8809 914 8843 948
rect 8877 914 8911 948
rect 8945 914 8979 948
rect 9013 914 9047 948
rect 9081 914 9115 948
rect 9149 914 9183 948
rect 9217 914 9251 948
rect 9285 914 9319 948
rect 9353 914 9365 948
rect 6365 903 9365 914
rect 65 818 3065 826
rect 65 784 95 818
rect 129 784 163 818
rect 197 784 231 818
rect 265 784 299 818
rect 333 784 367 818
rect 401 784 435 818
rect 469 784 503 818
rect 537 784 571 818
rect 605 784 639 818
rect 673 784 707 818
rect 741 784 775 818
rect 809 784 843 818
rect 877 784 911 818
rect 945 784 979 818
rect 1013 784 1047 818
rect 1081 784 1115 818
rect 1149 784 1183 818
rect 1217 784 1251 818
rect 1285 784 1319 818
rect 1353 784 1387 818
rect 1421 784 1455 818
rect 1489 784 1523 818
rect 1557 784 1591 818
rect 1625 784 1659 818
rect 1693 784 1727 818
rect 1761 784 1795 818
rect 1829 784 1863 818
rect 1897 784 1931 818
rect 1965 784 1999 818
rect 2033 784 2067 818
rect 2101 784 2135 818
rect 2169 784 2203 818
rect 2237 784 2271 818
rect 2305 784 2339 818
rect 2373 784 2407 818
rect 2441 784 2475 818
rect 2509 784 2543 818
rect 2577 784 2611 818
rect 2645 784 2679 818
rect 2713 784 2747 818
rect 2781 784 2815 818
rect 2849 784 2883 818
rect 2917 784 2951 818
rect 2985 784 3019 818
rect 3053 784 3065 818
rect 3215 818 6215 826
rect 65 773 3065 784
rect 3215 784 3245 818
rect 3279 784 3313 818
rect 3347 784 3381 818
rect 3415 784 3449 818
rect 3483 784 3517 818
rect 3551 784 3585 818
rect 3619 784 3653 818
rect 3687 784 3721 818
rect 3755 784 3789 818
rect 3823 784 3857 818
rect 3891 784 3925 818
rect 3959 784 3993 818
rect 4027 784 4061 818
rect 4095 784 4129 818
rect 4163 784 4197 818
rect 4231 784 4265 818
rect 4299 784 4333 818
rect 4367 784 4401 818
rect 4435 784 4469 818
rect 4503 784 4537 818
rect 4571 784 4605 818
rect 4639 784 4673 818
rect 4707 784 4741 818
rect 4775 784 4809 818
rect 4843 784 4877 818
rect 4911 784 4945 818
rect 4979 784 5013 818
rect 5047 784 5081 818
rect 5115 784 5149 818
rect 5183 784 5217 818
rect 5251 784 5285 818
rect 5319 784 5353 818
rect 5387 784 5421 818
rect 5455 784 5489 818
rect 5523 784 5557 818
rect 5591 784 5625 818
rect 5659 784 5693 818
rect 5727 784 5761 818
rect 5795 784 5829 818
rect 5863 784 5897 818
rect 5931 784 5965 818
rect 5999 784 6033 818
rect 6067 784 6101 818
rect 6135 784 6169 818
rect 6203 784 6215 818
rect 3215 773 6215 784
rect 9515 948 12515 959
rect 9515 914 9545 948
rect 9579 914 9613 948
rect 9647 914 9681 948
rect 9715 914 9749 948
rect 9783 914 9817 948
rect 9851 914 9885 948
rect 9919 914 9953 948
rect 9987 914 10021 948
rect 10055 914 10089 948
rect 10123 914 10157 948
rect 10191 914 10225 948
rect 10259 914 10293 948
rect 10327 914 10361 948
rect 10395 914 10429 948
rect 10463 914 10497 948
rect 10531 914 10565 948
rect 10599 914 10633 948
rect 10667 914 10701 948
rect 10735 914 10769 948
rect 10803 914 10837 948
rect 10871 914 10905 948
rect 10939 914 10973 948
rect 11007 914 11041 948
rect 11075 914 11109 948
rect 11143 914 11177 948
rect 11211 914 11245 948
rect 11279 914 11313 948
rect 11347 914 11381 948
rect 11415 914 11449 948
rect 11483 914 11517 948
rect 11551 914 11585 948
rect 11619 914 11653 948
rect 11687 914 11721 948
rect 11755 914 11789 948
rect 11823 914 11857 948
rect 11891 914 11925 948
rect 11959 914 11993 948
rect 12027 914 12061 948
rect 12095 914 12129 948
rect 12163 914 12197 948
rect 12231 914 12265 948
rect 12299 914 12333 948
rect 12367 914 12401 948
rect 12435 914 12469 948
rect 12503 914 12515 948
rect 9515 903 12515 914
rect 12665 948 15665 959
rect 12665 914 12695 948
rect 12729 914 12763 948
rect 12797 914 12831 948
rect 12865 914 12899 948
rect 12933 914 12967 948
rect 13001 914 13035 948
rect 13069 914 13103 948
rect 13137 914 13171 948
rect 13205 914 13239 948
rect 13273 914 13307 948
rect 13341 914 13375 948
rect 13409 914 13443 948
rect 13477 914 13511 948
rect 13545 914 13579 948
rect 13613 914 13647 948
rect 13681 914 13715 948
rect 13749 914 13783 948
rect 13817 914 13851 948
rect 13885 914 13919 948
rect 13953 914 13987 948
rect 14021 914 14055 948
rect 14089 914 14123 948
rect 14157 914 14191 948
rect 14225 914 14259 948
rect 14293 914 14327 948
rect 14361 914 14395 948
rect 14429 914 14463 948
rect 14497 914 14531 948
rect 14565 914 14599 948
rect 14633 914 14667 948
rect 14701 914 14735 948
rect 14769 914 14803 948
rect 14837 914 14871 948
rect 14905 914 14939 948
rect 14973 914 15007 948
rect 15041 914 15075 948
rect 15109 914 15143 948
rect 15177 914 15211 948
rect 15245 914 15279 948
rect 15313 914 15347 948
rect 15381 914 15415 948
rect 15449 914 15483 948
rect 15517 914 15551 948
rect 15585 914 15619 948
rect 15653 914 15665 948
rect 12665 903 15665 914
rect 15815 948 18815 959
rect 15815 914 15845 948
rect 15879 914 15913 948
rect 15947 914 15981 948
rect 16015 914 16049 948
rect 16083 914 16117 948
rect 16151 914 16185 948
rect 16219 914 16253 948
rect 16287 914 16321 948
rect 16355 914 16389 948
rect 16423 914 16457 948
rect 16491 914 16525 948
rect 16559 914 16593 948
rect 16627 914 16661 948
rect 16695 914 16729 948
rect 16763 914 16797 948
rect 16831 914 16865 948
rect 16899 914 16933 948
rect 16967 914 17001 948
rect 17035 914 17069 948
rect 17103 914 17137 948
rect 17171 914 17205 948
rect 17239 914 17273 948
rect 17307 914 17341 948
rect 17375 914 17409 948
rect 17443 914 17477 948
rect 17511 914 17545 948
rect 17579 914 17613 948
rect 17647 914 17681 948
rect 17715 914 17749 948
rect 17783 914 17817 948
rect 17851 914 17885 948
rect 17919 914 17953 948
rect 17987 914 18021 948
rect 18055 914 18089 948
rect 18123 914 18157 948
rect 18191 914 18225 948
rect 18259 914 18293 948
rect 18327 914 18361 948
rect 18395 914 18429 948
rect 18463 914 18497 948
rect 18531 914 18565 948
rect 18599 914 18633 948
rect 18667 914 18701 948
rect 18735 914 18769 948
rect 18803 914 18815 948
rect 15815 903 18815 914
rect 18965 948 21965 959
rect 18965 914 18995 948
rect 19029 914 19063 948
rect 19097 914 19131 948
rect 19165 914 19199 948
rect 19233 914 19267 948
rect 19301 914 19335 948
rect 19369 914 19403 948
rect 19437 914 19471 948
rect 19505 914 19539 948
rect 19573 914 19607 948
rect 19641 914 19675 948
rect 19709 914 19743 948
rect 19777 914 19811 948
rect 19845 914 19879 948
rect 19913 914 19947 948
rect 19981 914 20015 948
rect 20049 914 20083 948
rect 20117 914 20151 948
rect 20185 914 20219 948
rect 20253 914 20287 948
rect 20321 914 20355 948
rect 20389 914 20423 948
rect 20457 914 20491 948
rect 20525 914 20559 948
rect 20593 914 20627 948
rect 20661 914 20695 948
rect 20729 914 20763 948
rect 20797 914 20831 948
rect 20865 914 20899 948
rect 20933 914 20967 948
rect 21001 914 21035 948
rect 21069 914 21103 948
rect 21137 914 21171 948
rect 21205 914 21239 948
rect 21273 914 21307 948
rect 21341 914 21375 948
rect 21409 914 21443 948
rect 21477 914 21511 948
rect 21545 914 21579 948
rect 21613 914 21647 948
rect 21681 914 21715 948
rect 21749 914 21783 948
rect 21817 914 21851 948
rect 21885 914 21919 948
rect 21953 914 21965 948
rect 18965 903 21965 914
rect 6365 792 9365 803
rect 6365 758 6395 792
rect 6429 758 6463 792
rect 6497 758 6531 792
rect 6565 758 6599 792
rect 6633 758 6667 792
rect 6701 758 6735 792
rect 6769 758 6803 792
rect 6837 758 6871 792
rect 6905 758 6939 792
rect 6973 758 7007 792
rect 7041 758 7075 792
rect 7109 758 7143 792
rect 7177 758 7211 792
rect 7245 758 7279 792
rect 7313 758 7347 792
rect 7381 758 7415 792
rect 7449 758 7483 792
rect 7517 758 7551 792
rect 7585 758 7619 792
rect 7653 758 7687 792
rect 7721 758 7755 792
rect 7789 758 7823 792
rect 7857 758 7891 792
rect 7925 758 7959 792
rect 7993 758 8027 792
rect 8061 758 8095 792
rect 8129 758 8163 792
rect 8197 758 8231 792
rect 8265 758 8299 792
rect 8333 758 8367 792
rect 8401 758 8435 792
rect 8469 758 8503 792
rect 8537 758 8571 792
rect 8605 758 8639 792
rect 8673 758 8707 792
rect 8741 758 8775 792
rect 8809 758 8843 792
rect 8877 758 8911 792
rect 8945 758 8979 792
rect 9013 758 9047 792
rect 9081 758 9115 792
rect 9149 758 9183 792
rect 9217 758 9251 792
rect 9285 758 9319 792
rect 9353 758 9365 792
rect 6365 747 9365 758
rect 65 662 3065 673
rect 65 628 95 662
rect 129 628 163 662
rect 197 628 231 662
rect 265 628 299 662
rect 333 628 367 662
rect 401 628 435 662
rect 469 628 503 662
rect 537 628 571 662
rect 605 628 639 662
rect 673 628 707 662
rect 741 628 775 662
rect 809 628 843 662
rect 877 628 911 662
rect 945 628 979 662
rect 1013 628 1047 662
rect 1081 628 1115 662
rect 1149 628 1183 662
rect 1217 628 1251 662
rect 1285 628 1319 662
rect 1353 628 1387 662
rect 1421 628 1455 662
rect 1489 628 1523 662
rect 1557 628 1591 662
rect 1625 628 1659 662
rect 1693 628 1727 662
rect 1761 628 1795 662
rect 1829 628 1863 662
rect 1897 628 1931 662
rect 1965 628 1999 662
rect 2033 628 2067 662
rect 2101 628 2135 662
rect 2169 628 2203 662
rect 2237 628 2271 662
rect 2305 628 2339 662
rect 2373 628 2407 662
rect 2441 628 2475 662
rect 2509 628 2543 662
rect 2577 628 2611 662
rect 2645 628 2679 662
rect 2713 628 2747 662
rect 2781 628 2815 662
rect 2849 628 2883 662
rect 2917 628 2951 662
rect 2985 628 3019 662
rect 3053 628 3065 662
rect 65 620 3065 628
rect 3215 662 6215 673
rect 3215 628 3245 662
rect 3279 628 3313 662
rect 3347 628 3381 662
rect 3415 628 3449 662
rect 3483 628 3517 662
rect 3551 628 3585 662
rect 3619 628 3653 662
rect 3687 628 3721 662
rect 3755 628 3789 662
rect 3823 628 3857 662
rect 3891 628 3925 662
rect 3959 628 3993 662
rect 4027 628 4061 662
rect 4095 628 4129 662
rect 4163 628 4197 662
rect 4231 628 4265 662
rect 4299 628 4333 662
rect 4367 628 4401 662
rect 4435 628 4469 662
rect 4503 628 4537 662
rect 4571 628 4605 662
rect 4639 628 4673 662
rect 4707 628 4741 662
rect 4775 628 4809 662
rect 4843 628 4877 662
rect 4911 628 4945 662
rect 4979 628 5013 662
rect 5047 628 5081 662
rect 5115 628 5149 662
rect 5183 628 5217 662
rect 5251 628 5285 662
rect 5319 628 5353 662
rect 5387 628 5421 662
rect 5455 628 5489 662
rect 5523 628 5557 662
rect 5591 628 5625 662
rect 5659 628 5693 662
rect 5727 628 5761 662
rect 5795 628 5829 662
rect 5863 628 5897 662
rect 5931 628 5965 662
rect 5999 628 6033 662
rect 6067 628 6101 662
rect 6135 628 6169 662
rect 6203 628 6215 662
rect 9515 792 12515 803
rect 9515 758 9545 792
rect 9579 758 9613 792
rect 9647 758 9681 792
rect 9715 758 9749 792
rect 9783 758 9817 792
rect 9851 758 9885 792
rect 9919 758 9953 792
rect 9987 758 10021 792
rect 10055 758 10089 792
rect 10123 758 10157 792
rect 10191 758 10225 792
rect 10259 758 10293 792
rect 10327 758 10361 792
rect 10395 758 10429 792
rect 10463 758 10497 792
rect 10531 758 10565 792
rect 10599 758 10633 792
rect 10667 758 10701 792
rect 10735 758 10769 792
rect 10803 758 10837 792
rect 10871 758 10905 792
rect 10939 758 10973 792
rect 11007 758 11041 792
rect 11075 758 11109 792
rect 11143 758 11177 792
rect 11211 758 11245 792
rect 11279 758 11313 792
rect 11347 758 11381 792
rect 11415 758 11449 792
rect 11483 758 11517 792
rect 11551 758 11585 792
rect 11619 758 11653 792
rect 11687 758 11721 792
rect 11755 758 11789 792
rect 11823 758 11857 792
rect 11891 758 11925 792
rect 11959 758 11993 792
rect 12027 758 12061 792
rect 12095 758 12129 792
rect 12163 758 12197 792
rect 12231 758 12265 792
rect 12299 758 12333 792
rect 12367 758 12401 792
rect 12435 758 12469 792
rect 12503 758 12515 792
rect 9515 747 12515 758
rect 12665 792 15665 803
rect 12665 758 12695 792
rect 12729 758 12763 792
rect 12797 758 12831 792
rect 12865 758 12899 792
rect 12933 758 12967 792
rect 13001 758 13035 792
rect 13069 758 13103 792
rect 13137 758 13171 792
rect 13205 758 13239 792
rect 13273 758 13307 792
rect 13341 758 13375 792
rect 13409 758 13443 792
rect 13477 758 13511 792
rect 13545 758 13579 792
rect 13613 758 13647 792
rect 13681 758 13715 792
rect 13749 758 13783 792
rect 13817 758 13851 792
rect 13885 758 13919 792
rect 13953 758 13987 792
rect 14021 758 14055 792
rect 14089 758 14123 792
rect 14157 758 14191 792
rect 14225 758 14259 792
rect 14293 758 14327 792
rect 14361 758 14395 792
rect 14429 758 14463 792
rect 14497 758 14531 792
rect 14565 758 14599 792
rect 14633 758 14667 792
rect 14701 758 14735 792
rect 14769 758 14803 792
rect 14837 758 14871 792
rect 14905 758 14939 792
rect 14973 758 15007 792
rect 15041 758 15075 792
rect 15109 758 15143 792
rect 15177 758 15211 792
rect 15245 758 15279 792
rect 15313 758 15347 792
rect 15381 758 15415 792
rect 15449 758 15483 792
rect 15517 758 15551 792
rect 15585 758 15619 792
rect 15653 758 15665 792
rect 12665 747 15665 758
rect 15815 792 18815 803
rect 15815 758 15845 792
rect 15879 758 15913 792
rect 15947 758 15981 792
rect 16015 758 16049 792
rect 16083 758 16117 792
rect 16151 758 16185 792
rect 16219 758 16253 792
rect 16287 758 16321 792
rect 16355 758 16389 792
rect 16423 758 16457 792
rect 16491 758 16525 792
rect 16559 758 16593 792
rect 16627 758 16661 792
rect 16695 758 16729 792
rect 16763 758 16797 792
rect 16831 758 16865 792
rect 16899 758 16933 792
rect 16967 758 17001 792
rect 17035 758 17069 792
rect 17103 758 17137 792
rect 17171 758 17205 792
rect 17239 758 17273 792
rect 17307 758 17341 792
rect 17375 758 17409 792
rect 17443 758 17477 792
rect 17511 758 17545 792
rect 17579 758 17613 792
rect 17647 758 17681 792
rect 17715 758 17749 792
rect 17783 758 17817 792
rect 17851 758 17885 792
rect 17919 758 17953 792
rect 17987 758 18021 792
rect 18055 758 18089 792
rect 18123 758 18157 792
rect 18191 758 18225 792
rect 18259 758 18293 792
rect 18327 758 18361 792
rect 18395 758 18429 792
rect 18463 758 18497 792
rect 18531 758 18565 792
rect 18599 758 18633 792
rect 18667 758 18701 792
rect 18735 758 18769 792
rect 18803 758 18815 792
rect 15815 747 18815 758
rect 18965 792 21965 803
rect 18965 758 18995 792
rect 19029 758 19063 792
rect 19097 758 19131 792
rect 19165 758 19199 792
rect 19233 758 19267 792
rect 19301 758 19335 792
rect 19369 758 19403 792
rect 19437 758 19471 792
rect 19505 758 19539 792
rect 19573 758 19607 792
rect 19641 758 19675 792
rect 19709 758 19743 792
rect 19777 758 19811 792
rect 19845 758 19879 792
rect 19913 758 19947 792
rect 19981 758 20015 792
rect 20049 758 20083 792
rect 20117 758 20151 792
rect 20185 758 20219 792
rect 20253 758 20287 792
rect 20321 758 20355 792
rect 20389 758 20423 792
rect 20457 758 20491 792
rect 20525 758 20559 792
rect 20593 758 20627 792
rect 20661 758 20695 792
rect 20729 758 20763 792
rect 20797 758 20831 792
rect 20865 758 20899 792
rect 20933 758 20967 792
rect 21001 758 21035 792
rect 21069 758 21103 792
rect 21137 758 21171 792
rect 21205 758 21239 792
rect 21273 758 21307 792
rect 21341 758 21375 792
rect 21409 758 21443 792
rect 21477 758 21511 792
rect 21545 758 21579 792
rect 21613 758 21647 792
rect 21681 758 21715 792
rect 21749 758 21783 792
rect 21817 758 21851 792
rect 21885 758 21919 792
rect 21953 758 21965 792
rect 18965 747 21965 758
rect 22340 1170 24340 1181
rect 22340 1136 22390 1170
rect 22424 1136 22458 1170
rect 22492 1136 22526 1170
rect 22560 1136 22594 1170
rect 22628 1136 22662 1170
rect 22696 1136 22730 1170
rect 22764 1136 22798 1170
rect 22832 1136 22866 1170
rect 22900 1136 22934 1170
rect 22968 1136 23002 1170
rect 23036 1136 23070 1170
rect 23104 1136 23138 1170
rect 23172 1136 23206 1170
rect 23240 1136 23274 1170
rect 23308 1136 23342 1170
rect 23376 1136 23410 1170
rect 23444 1136 23478 1170
rect 23512 1136 23546 1170
rect 23580 1136 23614 1170
rect 23648 1136 23682 1170
rect 23716 1136 23750 1170
rect 23784 1136 23818 1170
rect 23852 1136 23886 1170
rect 23920 1136 23954 1170
rect 23988 1136 24022 1170
rect 24056 1136 24090 1170
rect 24124 1136 24158 1170
rect 24192 1136 24226 1170
rect 24260 1136 24294 1170
rect 24328 1136 24340 1170
rect 22340 1125 24340 1136
rect 22340 1014 24340 1025
rect 22340 980 22390 1014
rect 22424 980 22458 1014
rect 22492 980 22526 1014
rect 22560 980 22594 1014
rect 22628 980 22662 1014
rect 22696 980 22730 1014
rect 22764 980 22798 1014
rect 22832 980 22866 1014
rect 22900 980 22934 1014
rect 22968 980 23002 1014
rect 23036 980 23070 1014
rect 23104 980 23138 1014
rect 23172 980 23206 1014
rect 23240 980 23274 1014
rect 23308 980 23342 1014
rect 23376 980 23410 1014
rect 23444 980 23478 1014
rect 23512 980 23546 1014
rect 23580 980 23614 1014
rect 23648 980 23682 1014
rect 23716 980 23750 1014
rect 23784 980 23818 1014
rect 23852 980 23886 1014
rect 23920 980 23954 1014
rect 23988 980 24022 1014
rect 24056 980 24090 1014
rect 24124 980 24158 1014
rect 24192 980 24226 1014
rect 24260 980 24294 1014
rect 24328 980 24340 1014
rect 22340 969 24340 980
rect 22340 858 24340 869
rect 22340 824 22390 858
rect 22424 824 22458 858
rect 22492 824 22526 858
rect 22560 824 22594 858
rect 22628 824 22662 858
rect 22696 824 22730 858
rect 22764 824 22798 858
rect 22832 824 22866 858
rect 22900 824 22934 858
rect 22968 824 23002 858
rect 23036 824 23070 858
rect 23104 824 23138 858
rect 23172 824 23206 858
rect 23240 824 23274 858
rect 23308 824 23342 858
rect 23376 824 23410 858
rect 23444 824 23478 858
rect 23512 824 23546 858
rect 23580 824 23614 858
rect 23648 824 23682 858
rect 23716 824 23750 858
rect 23784 824 23818 858
rect 23852 824 23886 858
rect 23920 824 23954 858
rect 23988 824 24022 858
rect 24056 824 24090 858
rect 24124 824 24158 858
rect 24192 824 24226 858
rect 24260 824 24294 858
rect 24328 824 24340 858
rect 22340 813 24340 824
rect 22340 702 24340 713
rect 22340 668 22390 702
rect 22424 668 22458 702
rect 22492 668 22526 702
rect 22560 668 22594 702
rect 22628 668 22662 702
rect 22696 668 22730 702
rect 22764 668 22798 702
rect 22832 668 22866 702
rect 22900 668 22934 702
rect 22968 668 23002 702
rect 23036 668 23070 702
rect 23104 668 23138 702
rect 23172 668 23206 702
rect 23240 668 23274 702
rect 23308 668 23342 702
rect 23376 668 23410 702
rect 23444 668 23478 702
rect 23512 668 23546 702
rect 23580 668 23614 702
rect 23648 668 23682 702
rect 23716 668 23750 702
rect 23784 668 23818 702
rect 23852 668 23886 702
rect 23920 668 23954 702
rect 23988 668 24022 702
rect 24056 668 24090 702
rect 24124 668 24158 702
rect 24192 668 24226 702
rect 24260 668 24294 702
rect 24328 668 24340 702
rect 22340 660 24340 668
rect 3215 620 6215 628
rect 6365 636 9365 647
rect 6365 602 6395 636
rect 6429 602 6463 636
rect 6497 602 6531 636
rect 6565 602 6599 636
rect 6633 602 6667 636
rect 6701 602 6735 636
rect 6769 602 6803 636
rect 6837 602 6871 636
rect 6905 602 6939 636
rect 6973 602 7007 636
rect 7041 602 7075 636
rect 7109 602 7143 636
rect 7177 602 7211 636
rect 7245 602 7279 636
rect 7313 602 7347 636
rect 7381 602 7415 636
rect 7449 602 7483 636
rect 7517 602 7551 636
rect 7585 602 7619 636
rect 7653 602 7687 636
rect 7721 602 7755 636
rect 7789 602 7823 636
rect 7857 602 7891 636
rect 7925 602 7959 636
rect 7993 602 8027 636
rect 8061 602 8095 636
rect 8129 602 8163 636
rect 8197 602 8231 636
rect 8265 602 8299 636
rect 8333 602 8367 636
rect 8401 602 8435 636
rect 8469 602 8503 636
rect 8537 602 8571 636
rect 8605 602 8639 636
rect 8673 602 8707 636
rect 8741 602 8775 636
rect 8809 602 8843 636
rect 8877 602 8911 636
rect 8945 602 8979 636
rect 9013 602 9047 636
rect 9081 602 9115 636
rect 9149 602 9183 636
rect 9217 602 9251 636
rect 9285 602 9319 636
rect 9353 602 9365 636
rect 6365 594 9365 602
rect 9515 636 12515 647
rect 9515 602 9545 636
rect 9579 602 9613 636
rect 9647 602 9681 636
rect 9715 602 9749 636
rect 9783 602 9817 636
rect 9851 602 9885 636
rect 9919 602 9953 636
rect 9987 602 10021 636
rect 10055 602 10089 636
rect 10123 602 10157 636
rect 10191 602 10225 636
rect 10259 602 10293 636
rect 10327 602 10361 636
rect 10395 602 10429 636
rect 10463 602 10497 636
rect 10531 602 10565 636
rect 10599 602 10633 636
rect 10667 602 10701 636
rect 10735 602 10769 636
rect 10803 602 10837 636
rect 10871 602 10905 636
rect 10939 602 10973 636
rect 11007 602 11041 636
rect 11075 602 11109 636
rect 11143 602 11177 636
rect 11211 602 11245 636
rect 11279 602 11313 636
rect 11347 602 11381 636
rect 11415 602 11449 636
rect 11483 602 11517 636
rect 11551 602 11585 636
rect 11619 602 11653 636
rect 11687 602 11721 636
rect 11755 602 11789 636
rect 11823 602 11857 636
rect 11891 602 11925 636
rect 11959 602 11993 636
rect 12027 602 12061 636
rect 12095 602 12129 636
rect 12163 602 12197 636
rect 12231 602 12265 636
rect 12299 602 12333 636
rect 12367 602 12401 636
rect 12435 602 12469 636
rect 12503 602 12515 636
rect 9515 594 12515 602
rect 12665 636 15665 647
rect 12665 602 12695 636
rect 12729 602 12763 636
rect 12797 602 12831 636
rect 12865 602 12899 636
rect 12933 602 12967 636
rect 13001 602 13035 636
rect 13069 602 13103 636
rect 13137 602 13171 636
rect 13205 602 13239 636
rect 13273 602 13307 636
rect 13341 602 13375 636
rect 13409 602 13443 636
rect 13477 602 13511 636
rect 13545 602 13579 636
rect 13613 602 13647 636
rect 13681 602 13715 636
rect 13749 602 13783 636
rect 13817 602 13851 636
rect 13885 602 13919 636
rect 13953 602 13987 636
rect 14021 602 14055 636
rect 14089 602 14123 636
rect 14157 602 14191 636
rect 14225 602 14259 636
rect 14293 602 14327 636
rect 14361 602 14395 636
rect 14429 602 14463 636
rect 14497 602 14531 636
rect 14565 602 14599 636
rect 14633 602 14667 636
rect 14701 602 14735 636
rect 14769 602 14803 636
rect 14837 602 14871 636
rect 14905 602 14939 636
rect 14973 602 15007 636
rect 15041 602 15075 636
rect 15109 602 15143 636
rect 15177 602 15211 636
rect 15245 602 15279 636
rect 15313 602 15347 636
rect 15381 602 15415 636
rect 15449 602 15483 636
rect 15517 602 15551 636
rect 15585 602 15619 636
rect 15653 602 15665 636
rect 12665 594 15665 602
rect 15815 636 18815 647
rect 15815 602 15845 636
rect 15879 602 15913 636
rect 15947 602 15981 636
rect 16015 602 16049 636
rect 16083 602 16117 636
rect 16151 602 16185 636
rect 16219 602 16253 636
rect 16287 602 16321 636
rect 16355 602 16389 636
rect 16423 602 16457 636
rect 16491 602 16525 636
rect 16559 602 16593 636
rect 16627 602 16661 636
rect 16695 602 16729 636
rect 16763 602 16797 636
rect 16831 602 16865 636
rect 16899 602 16933 636
rect 16967 602 17001 636
rect 17035 602 17069 636
rect 17103 602 17137 636
rect 17171 602 17205 636
rect 17239 602 17273 636
rect 17307 602 17341 636
rect 17375 602 17409 636
rect 17443 602 17477 636
rect 17511 602 17545 636
rect 17579 602 17613 636
rect 17647 602 17681 636
rect 17715 602 17749 636
rect 17783 602 17817 636
rect 17851 602 17885 636
rect 17919 602 17953 636
rect 17987 602 18021 636
rect 18055 602 18089 636
rect 18123 602 18157 636
rect 18191 602 18225 636
rect 18259 602 18293 636
rect 18327 602 18361 636
rect 18395 602 18429 636
rect 18463 602 18497 636
rect 18531 602 18565 636
rect 18599 602 18633 636
rect 18667 602 18701 636
rect 18735 602 18769 636
rect 18803 602 18815 636
rect 15815 594 18815 602
rect 18965 636 21965 647
rect 18965 602 18995 636
rect 19029 602 19063 636
rect 19097 602 19131 636
rect 19165 602 19199 636
rect 19233 602 19267 636
rect 19301 602 19335 636
rect 19369 602 19403 636
rect 19437 602 19471 636
rect 19505 602 19539 636
rect 19573 602 19607 636
rect 19641 602 19675 636
rect 19709 602 19743 636
rect 19777 602 19811 636
rect 19845 602 19879 636
rect 19913 602 19947 636
rect 19981 602 20015 636
rect 20049 602 20083 636
rect 20117 602 20151 636
rect 20185 602 20219 636
rect 20253 602 20287 636
rect 20321 602 20355 636
rect 20389 602 20423 636
rect 20457 602 20491 636
rect 20525 602 20559 636
rect 20593 602 20627 636
rect 20661 602 20695 636
rect 20729 602 20763 636
rect 20797 602 20831 636
rect 20865 602 20899 636
rect 20933 602 20967 636
rect 21001 602 21035 636
rect 21069 602 21103 636
rect 21137 602 21171 636
rect 21205 602 21239 636
rect 21273 602 21307 636
rect 21341 602 21375 636
rect 21409 602 21443 636
rect 21477 602 21511 636
rect 21545 602 21579 636
rect 21613 602 21647 636
rect 21681 602 21715 636
rect 21749 602 21783 636
rect 21817 602 21851 636
rect 21885 602 21919 636
rect 21953 602 21965 636
rect 18965 594 21965 602
<< mvpdiffc >>
rect 22390 2072 22424 2106
rect 22458 2072 22492 2106
rect 22526 2072 22560 2106
rect 22594 2072 22628 2106
rect 22662 2072 22696 2106
rect 22730 2072 22764 2106
rect 22798 2072 22832 2106
rect 22866 2072 22900 2106
rect 22934 2072 22968 2106
rect 23002 2072 23036 2106
rect 23070 2072 23104 2106
rect 23138 2072 23172 2106
rect 23206 2072 23240 2106
rect 23274 2072 23308 2106
rect 23342 2072 23376 2106
rect 23410 2072 23444 2106
rect 23478 2072 23512 2106
rect 23546 2072 23580 2106
rect 23614 2072 23648 2106
rect 23682 2072 23716 2106
rect 23750 2072 23784 2106
rect 23818 2072 23852 2106
rect 23886 2072 23920 2106
rect 23954 2072 23988 2106
rect 24022 2072 24056 2106
rect 24090 2072 24124 2106
rect 24158 2072 24192 2106
rect 24226 2072 24260 2106
rect 24294 2072 24328 2106
rect 22390 1916 22424 1950
rect 22458 1916 22492 1950
rect 22526 1916 22560 1950
rect 22594 1916 22628 1950
rect 22662 1916 22696 1950
rect 22730 1916 22764 1950
rect 22798 1916 22832 1950
rect 22866 1916 22900 1950
rect 22934 1916 22968 1950
rect 23002 1916 23036 1950
rect 23070 1916 23104 1950
rect 23138 1916 23172 1950
rect 23206 1916 23240 1950
rect 23274 1916 23308 1950
rect 23342 1916 23376 1950
rect 23410 1916 23444 1950
rect 23478 1916 23512 1950
rect 23546 1916 23580 1950
rect 23614 1916 23648 1950
rect 23682 1916 23716 1950
rect 23750 1916 23784 1950
rect 23818 1916 23852 1950
rect 23886 1916 23920 1950
rect 23954 1916 23988 1950
rect 24022 1916 24056 1950
rect 24090 1916 24124 1950
rect 24158 1916 24192 1950
rect 24226 1916 24260 1950
rect 24294 1916 24328 1950
rect 22390 1760 22424 1794
rect 22458 1760 22492 1794
rect 22526 1760 22560 1794
rect 22594 1760 22628 1794
rect 22662 1760 22696 1794
rect 22730 1760 22764 1794
rect 22798 1760 22832 1794
rect 22866 1760 22900 1794
rect 22934 1760 22968 1794
rect 23002 1760 23036 1794
rect 23070 1760 23104 1794
rect 23138 1760 23172 1794
rect 23206 1760 23240 1794
rect 23274 1760 23308 1794
rect 23342 1760 23376 1794
rect 23410 1760 23444 1794
rect 23478 1760 23512 1794
rect 23546 1760 23580 1794
rect 23614 1760 23648 1794
rect 23682 1760 23716 1794
rect 23750 1760 23784 1794
rect 23818 1760 23852 1794
rect 23886 1760 23920 1794
rect 23954 1760 23988 1794
rect 24022 1760 24056 1794
rect 24090 1760 24124 1794
rect 24158 1760 24192 1794
rect 24226 1760 24260 1794
rect 24294 1760 24328 1794
rect 22390 1604 22424 1638
rect 22458 1604 22492 1638
rect 22526 1604 22560 1638
rect 22594 1604 22628 1638
rect 22662 1604 22696 1638
rect 22730 1604 22764 1638
rect 22798 1604 22832 1638
rect 22866 1604 22900 1638
rect 22934 1604 22968 1638
rect 23002 1604 23036 1638
rect 23070 1604 23104 1638
rect 23138 1604 23172 1638
rect 23206 1604 23240 1638
rect 23274 1604 23308 1638
rect 23342 1604 23376 1638
rect 23410 1604 23444 1638
rect 23478 1604 23512 1638
rect 23546 1604 23580 1638
rect 23614 1604 23648 1638
rect 23682 1604 23716 1638
rect 23750 1604 23784 1638
rect 23818 1604 23852 1638
rect 23886 1604 23920 1638
rect 23954 1604 23988 1638
rect 24022 1604 24056 1638
rect 24090 1604 24124 1638
rect 24158 1604 24192 1638
rect 24226 1604 24260 1638
rect 24294 1604 24328 1638
rect 22390 1448 22424 1482
rect 22458 1448 22492 1482
rect 22526 1448 22560 1482
rect 22594 1448 22628 1482
rect 22662 1448 22696 1482
rect 22730 1448 22764 1482
rect 22798 1448 22832 1482
rect 22866 1448 22900 1482
rect 22934 1448 22968 1482
rect 23002 1448 23036 1482
rect 23070 1448 23104 1482
rect 23138 1448 23172 1482
rect 23206 1448 23240 1482
rect 23274 1448 23308 1482
rect 23342 1448 23376 1482
rect 23410 1448 23444 1482
rect 23478 1448 23512 1482
rect 23546 1448 23580 1482
rect 23614 1448 23648 1482
rect 23682 1448 23716 1482
rect 23750 1448 23784 1482
rect 23818 1448 23852 1482
rect 23886 1448 23920 1482
rect 23954 1448 23988 1482
rect 24022 1448 24056 1482
rect 24090 1448 24124 1482
rect 24158 1448 24192 1482
rect 24226 1448 24260 1482
rect 24294 1448 24328 1482
rect 22390 1292 22424 1326
rect 22458 1292 22492 1326
rect 22526 1292 22560 1326
rect 22594 1292 22628 1326
rect 22662 1292 22696 1326
rect 22730 1292 22764 1326
rect 22798 1292 22832 1326
rect 22866 1292 22900 1326
rect 22934 1292 22968 1326
rect 23002 1292 23036 1326
rect 23070 1292 23104 1326
rect 23138 1292 23172 1326
rect 23206 1292 23240 1326
rect 23274 1292 23308 1326
rect 23342 1292 23376 1326
rect 23410 1292 23444 1326
rect 23478 1292 23512 1326
rect 23546 1292 23580 1326
rect 23614 1292 23648 1326
rect 23682 1292 23716 1326
rect 23750 1292 23784 1326
rect 23818 1292 23852 1326
rect 23886 1292 23920 1326
rect 23954 1292 23988 1326
rect 24022 1292 24056 1326
rect 24090 1292 24124 1326
rect 24158 1292 24192 1326
rect 24226 1292 24260 1326
rect 24294 1292 24328 1326
rect 6395 1226 6429 1260
rect 6463 1226 6497 1260
rect 6531 1226 6565 1260
rect 6599 1226 6633 1260
rect 6667 1226 6701 1260
rect 6735 1226 6769 1260
rect 6803 1226 6837 1260
rect 6871 1226 6905 1260
rect 6939 1226 6973 1260
rect 7007 1226 7041 1260
rect 7075 1226 7109 1260
rect 7143 1226 7177 1260
rect 7211 1226 7245 1260
rect 7279 1226 7313 1260
rect 7347 1226 7381 1260
rect 7415 1226 7449 1260
rect 7483 1226 7517 1260
rect 7551 1226 7585 1260
rect 7619 1226 7653 1260
rect 7687 1226 7721 1260
rect 7755 1226 7789 1260
rect 7823 1226 7857 1260
rect 7891 1226 7925 1260
rect 7959 1226 7993 1260
rect 8027 1226 8061 1260
rect 8095 1226 8129 1260
rect 8163 1226 8197 1260
rect 8231 1226 8265 1260
rect 8299 1226 8333 1260
rect 8367 1226 8401 1260
rect 8435 1226 8469 1260
rect 8503 1226 8537 1260
rect 8571 1226 8605 1260
rect 8639 1226 8673 1260
rect 8707 1226 8741 1260
rect 8775 1226 8809 1260
rect 8843 1226 8877 1260
rect 8911 1226 8945 1260
rect 8979 1226 9013 1260
rect 9047 1226 9081 1260
rect 9115 1226 9149 1260
rect 9183 1226 9217 1260
rect 9251 1226 9285 1260
rect 9319 1226 9353 1260
rect 9545 1226 9579 1260
rect 9613 1226 9647 1260
rect 9681 1226 9715 1260
rect 9749 1226 9783 1260
rect 9817 1226 9851 1260
rect 9885 1226 9919 1260
rect 9953 1226 9987 1260
rect 10021 1226 10055 1260
rect 10089 1226 10123 1260
rect 10157 1226 10191 1260
rect 10225 1226 10259 1260
rect 10293 1226 10327 1260
rect 10361 1226 10395 1260
rect 10429 1226 10463 1260
rect 10497 1226 10531 1260
rect 10565 1226 10599 1260
rect 10633 1226 10667 1260
rect 10701 1226 10735 1260
rect 10769 1226 10803 1260
rect 10837 1226 10871 1260
rect 10905 1226 10939 1260
rect 10973 1226 11007 1260
rect 11041 1226 11075 1260
rect 11109 1226 11143 1260
rect 11177 1226 11211 1260
rect 11245 1226 11279 1260
rect 11313 1226 11347 1260
rect 11381 1226 11415 1260
rect 11449 1226 11483 1260
rect 11517 1226 11551 1260
rect 11585 1226 11619 1260
rect 11653 1226 11687 1260
rect 11721 1226 11755 1260
rect 11789 1226 11823 1260
rect 11857 1226 11891 1260
rect 11925 1226 11959 1260
rect 11993 1226 12027 1260
rect 12061 1226 12095 1260
rect 12129 1226 12163 1260
rect 12197 1226 12231 1260
rect 12265 1226 12299 1260
rect 12333 1226 12367 1260
rect 12401 1226 12435 1260
rect 12469 1226 12503 1260
rect 12695 1226 12729 1260
rect 12763 1226 12797 1260
rect 12831 1226 12865 1260
rect 12899 1226 12933 1260
rect 12967 1226 13001 1260
rect 13035 1226 13069 1260
rect 13103 1226 13137 1260
rect 13171 1226 13205 1260
rect 13239 1226 13273 1260
rect 13307 1226 13341 1260
rect 13375 1226 13409 1260
rect 13443 1226 13477 1260
rect 13511 1226 13545 1260
rect 13579 1226 13613 1260
rect 13647 1226 13681 1260
rect 13715 1226 13749 1260
rect 13783 1226 13817 1260
rect 13851 1226 13885 1260
rect 13919 1226 13953 1260
rect 13987 1226 14021 1260
rect 14055 1226 14089 1260
rect 14123 1226 14157 1260
rect 14191 1226 14225 1260
rect 14259 1226 14293 1260
rect 14327 1226 14361 1260
rect 14395 1226 14429 1260
rect 14463 1226 14497 1260
rect 14531 1226 14565 1260
rect 14599 1226 14633 1260
rect 14667 1226 14701 1260
rect 14735 1226 14769 1260
rect 14803 1226 14837 1260
rect 14871 1226 14905 1260
rect 14939 1226 14973 1260
rect 15007 1226 15041 1260
rect 15075 1226 15109 1260
rect 15143 1226 15177 1260
rect 15211 1226 15245 1260
rect 15279 1226 15313 1260
rect 15347 1226 15381 1260
rect 15415 1226 15449 1260
rect 15483 1226 15517 1260
rect 15551 1226 15585 1260
rect 15619 1226 15653 1260
rect 15845 1226 15879 1260
rect 15913 1226 15947 1260
rect 15981 1226 16015 1260
rect 16049 1226 16083 1260
rect 16117 1226 16151 1260
rect 16185 1226 16219 1260
rect 16253 1226 16287 1260
rect 16321 1226 16355 1260
rect 16389 1226 16423 1260
rect 16457 1226 16491 1260
rect 16525 1226 16559 1260
rect 16593 1226 16627 1260
rect 16661 1226 16695 1260
rect 16729 1226 16763 1260
rect 16797 1226 16831 1260
rect 16865 1226 16899 1260
rect 16933 1226 16967 1260
rect 17001 1226 17035 1260
rect 17069 1226 17103 1260
rect 17137 1226 17171 1260
rect 17205 1226 17239 1260
rect 17273 1226 17307 1260
rect 17341 1226 17375 1260
rect 17409 1226 17443 1260
rect 17477 1226 17511 1260
rect 17545 1226 17579 1260
rect 17613 1226 17647 1260
rect 17681 1226 17715 1260
rect 17749 1226 17783 1260
rect 17817 1226 17851 1260
rect 17885 1226 17919 1260
rect 17953 1226 17987 1260
rect 18021 1226 18055 1260
rect 18089 1226 18123 1260
rect 18157 1226 18191 1260
rect 18225 1226 18259 1260
rect 18293 1226 18327 1260
rect 18361 1226 18395 1260
rect 18429 1226 18463 1260
rect 18497 1226 18531 1260
rect 18565 1226 18599 1260
rect 18633 1226 18667 1260
rect 18701 1226 18735 1260
rect 18769 1226 18803 1260
rect 18995 1226 19029 1260
rect 19063 1226 19097 1260
rect 19131 1226 19165 1260
rect 19199 1226 19233 1260
rect 19267 1226 19301 1260
rect 19335 1226 19369 1260
rect 19403 1226 19437 1260
rect 19471 1226 19505 1260
rect 19539 1226 19573 1260
rect 19607 1226 19641 1260
rect 19675 1226 19709 1260
rect 19743 1226 19777 1260
rect 19811 1226 19845 1260
rect 19879 1226 19913 1260
rect 19947 1226 19981 1260
rect 20015 1226 20049 1260
rect 20083 1226 20117 1260
rect 20151 1226 20185 1260
rect 20219 1226 20253 1260
rect 20287 1226 20321 1260
rect 20355 1226 20389 1260
rect 20423 1226 20457 1260
rect 20491 1226 20525 1260
rect 20559 1226 20593 1260
rect 20627 1226 20661 1260
rect 20695 1226 20729 1260
rect 20763 1226 20797 1260
rect 20831 1226 20865 1260
rect 20899 1226 20933 1260
rect 20967 1226 21001 1260
rect 21035 1226 21069 1260
rect 21103 1226 21137 1260
rect 21171 1226 21205 1260
rect 21239 1226 21273 1260
rect 21307 1226 21341 1260
rect 21375 1226 21409 1260
rect 21443 1226 21477 1260
rect 21511 1226 21545 1260
rect 21579 1226 21613 1260
rect 21647 1226 21681 1260
rect 21715 1226 21749 1260
rect 21783 1226 21817 1260
rect 21851 1226 21885 1260
rect 21919 1226 21953 1260
rect 6395 1070 6429 1104
rect 6463 1070 6497 1104
rect 6531 1070 6565 1104
rect 6599 1070 6633 1104
rect 6667 1070 6701 1104
rect 6735 1070 6769 1104
rect 6803 1070 6837 1104
rect 6871 1070 6905 1104
rect 6939 1070 6973 1104
rect 7007 1070 7041 1104
rect 7075 1070 7109 1104
rect 7143 1070 7177 1104
rect 7211 1070 7245 1104
rect 7279 1070 7313 1104
rect 7347 1070 7381 1104
rect 7415 1070 7449 1104
rect 7483 1070 7517 1104
rect 7551 1070 7585 1104
rect 7619 1070 7653 1104
rect 7687 1070 7721 1104
rect 7755 1070 7789 1104
rect 7823 1070 7857 1104
rect 7891 1070 7925 1104
rect 7959 1070 7993 1104
rect 8027 1070 8061 1104
rect 8095 1070 8129 1104
rect 8163 1070 8197 1104
rect 8231 1070 8265 1104
rect 8299 1070 8333 1104
rect 8367 1070 8401 1104
rect 8435 1070 8469 1104
rect 8503 1070 8537 1104
rect 8571 1070 8605 1104
rect 8639 1070 8673 1104
rect 8707 1070 8741 1104
rect 8775 1070 8809 1104
rect 8843 1070 8877 1104
rect 8911 1070 8945 1104
rect 8979 1070 9013 1104
rect 9047 1070 9081 1104
rect 9115 1070 9149 1104
rect 9183 1070 9217 1104
rect 9251 1070 9285 1104
rect 9319 1070 9353 1104
rect 9545 1070 9579 1104
rect 9613 1070 9647 1104
rect 9681 1070 9715 1104
rect 9749 1070 9783 1104
rect 9817 1070 9851 1104
rect 9885 1070 9919 1104
rect 9953 1070 9987 1104
rect 10021 1070 10055 1104
rect 10089 1070 10123 1104
rect 10157 1070 10191 1104
rect 10225 1070 10259 1104
rect 10293 1070 10327 1104
rect 10361 1070 10395 1104
rect 10429 1070 10463 1104
rect 10497 1070 10531 1104
rect 10565 1070 10599 1104
rect 10633 1070 10667 1104
rect 10701 1070 10735 1104
rect 10769 1070 10803 1104
rect 10837 1070 10871 1104
rect 10905 1070 10939 1104
rect 10973 1070 11007 1104
rect 11041 1070 11075 1104
rect 11109 1070 11143 1104
rect 11177 1070 11211 1104
rect 11245 1070 11279 1104
rect 11313 1070 11347 1104
rect 11381 1070 11415 1104
rect 11449 1070 11483 1104
rect 11517 1070 11551 1104
rect 11585 1070 11619 1104
rect 11653 1070 11687 1104
rect 11721 1070 11755 1104
rect 11789 1070 11823 1104
rect 11857 1070 11891 1104
rect 11925 1070 11959 1104
rect 11993 1070 12027 1104
rect 12061 1070 12095 1104
rect 12129 1070 12163 1104
rect 12197 1070 12231 1104
rect 12265 1070 12299 1104
rect 12333 1070 12367 1104
rect 12401 1070 12435 1104
rect 12469 1070 12503 1104
rect 12695 1070 12729 1104
rect 12763 1070 12797 1104
rect 12831 1070 12865 1104
rect 12899 1070 12933 1104
rect 12967 1070 13001 1104
rect 13035 1070 13069 1104
rect 13103 1070 13137 1104
rect 13171 1070 13205 1104
rect 13239 1070 13273 1104
rect 13307 1070 13341 1104
rect 13375 1070 13409 1104
rect 13443 1070 13477 1104
rect 13511 1070 13545 1104
rect 13579 1070 13613 1104
rect 13647 1070 13681 1104
rect 13715 1070 13749 1104
rect 13783 1070 13817 1104
rect 13851 1070 13885 1104
rect 13919 1070 13953 1104
rect 13987 1070 14021 1104
rect 14055 1070 14089 1104
rect 14123 1070 14157 1104
rect 14191 1070 14225 1104
rect 14259 1070 14293 1104
rect 14327 1070 14361 1104
rect 14395 1070 14429 1104
rect 14463 1070 14497 1104
rect 14531 1070 14565 1104
rect 14599 1070 14633 1104
rect 14667 1070 14701 1104
rect 14735 1070 14769 1104
rect 14803 1070 14837 1104
rect 14871 1070 14905 1104
rect 14939 1070 14973 1104
rect 15007 1070 15041 1104
rect 15075 1070 15109 1104
rect 15143 1070 15177 1104
rect 15211 1070 15245 1104
rect 15279 1070 15313 1104
rect 15347 1070 15381 1104
rect 15415 1070 15449 1104
rect 15483 1070 15517 1104
rect 15551 1070 15585 1104
rect 15619 1070 15653 1104
rect 15845 1070 15879 1104
rect 15913 1070 15947 1104
rect 15981 1070 16015 1104
rect 16049 1070 16083 1104
rect 16117 1070 16151 1104
rect 16185 1070 16219 1104
rect 16253 1070 16287 1104
rect 16321 1070 16355 1104
rect 16389 1070 16423 1104
rect 16457 1070 16491 1104
rect 16525 1070 16559 1104
rect 16593 1070 16627 1104
rect 16661 1070 16695 1104
rect 16729 1070 16763 1104
rect 16797 1070 16831 1104
rect 16865 1070 16899 1104
rect 16933 1070 16967 1104
rect 17001 1070 17035 1104
rect 17069 1070 17103 1104
rect 17137 1070 17171 1104
rect 17205 1070 17239 1104
rect 17273 1070 17307 1104
rect 17341 1070 17375 1104
rect 17409 1070 17443 1104
rect 17477 1070 17511 1104
rect 17545 1070 17579 1104
rect 17613 1070 17647 1104
rect 17681 1070 17715 1104
rect 17749 1070 17783 1104
rect 17817 1070 17851 1104
rect 17885 1070 17919 1104
rect 17953 1070 17987 1104
rect 18021 1070 18055 1104
rect 18089 1070 18123 1104
rect 18157 1070 18191 1104
rect 18225 1070 18259 1104
rect 18293 1070 18327 1104
rect 18361 1070 18395 1104
rect 18429 1070 18463 1104
rect 18497 1070 18531 1104
rect 18565 1070 18599 1104
rect 18633 1070 18667 1104
rect 18701 1070 18735 1104
rect 18769 1070 18803 1104
rect 18995 1070 19029 1104
rect 19063 1070 19097 1104
rect 19131 1070 19165 1104
rect 19199 1070 19233 1104
rect 19267 1070 19301 1104
rect 19335 1070 19369 1104
rect 19403 1070 19437 1104
rect 19471 1070 19505 1104
rect 19539 1070 19573 1104
rect 19607 1070 19641 1104
rect 19675 1070 19709 1104
rect 19743 1070 19777 1104
rect 19811 1070 19845 1104
rect 19879 1070 19913 1104
rect 19947 1070 19981 1104
rect 20015 1070 20049 1104
rect 20083 1070 20117 1104
rect 20151 1070 20185 1104
rect 20219 1070 20253 1104
rect 20287 1070 20321 1104
rect 20355 1070 20389 1104
rect 20423 1070 20457 1104
rect 20491 1070 20525 1104
rect 20559 1070 20593 1104
rect 20627 1070 20661 1104
rect 20695 1070 20729 1104
rect 20763 1070 20797 1104
rect 20831 1070 20865 1104
rect 20899 1070 20933 1104
rect 20967 1070 21001 1104
rect 21035 1070 21069 1104
rect 21103 1070 21137 1104
rect 21171 1070 21205 1104
rect 21239 1070 21273 1104
rect 21307 1070 21341 1104
rect 21375 1070 21409 1104
rect 21443 1070 21477 1104
rect 21511 1070 21545 1104
rect 21579 1070 21613 1104
rect 21647 1070 21681 1104
rect 21715 1070 21749 1104
rect 21783 1070 21817 1104
rect 21851 1070 21885 1104
rect 21919 1070 21953 1104
rect 6395 914 6429 948
rect 6463 914 6497 948
rect 6531 914 6565 948
rect 6599 914 6633 948
rect 6667 914 6701 948
rect 6735 914 6769 948
rect 6803 914 6837 948
rect 6871 914 6905 948
rect 6939 914 6973 948
rect 7007 914 7041 948
rect 7075 914 7109 948
rect 7143 914 7177 948
rect 7211 914 7245 948
rect 7279 914 7313 948
rect 7347 914 7381 948
rect 7415 914 7449 948
rect 7483 914 7517 948
rect 7551 914 7585 948
rect 7619 914 7653 948
rect 7687 914 7721 948
rect 7755 914 7789 948
rect 7823 914 7857 948
rect 7891 914 7925 948
rect 7959 914 7993 948
rect 8027 914 8061 948
rect 8095 914 8129 948
rect 8163 914 8197 948
rect 8231 914 8265 948
rect 8299 914 8333 948
rect 8367 914 8401 948
rect 8435 914 8469 948
rect 8503 914 8537 948
rect 8571 914 8605 948
rect 8639 914 8673 948
rect 8707 914 8741 948
rect 8775 914 8809 948
rect 8843 914 8877 948
rect 8911 914 8945 948
rect 8979 914 9013 948
rect 9047 914 9081 948
rect 9115 914 9149 948
rect 9183 914 9217 948
rect 9251 914 9285 948
rect 9319 914 9353 948
rect 95 784 129 818
rect 163 784 197 818
rect 231 784 265 818
rect 299 784 333 818
rect 367 784 401 818
rect 435 784 469 818
rect 503 784 537 818
rect 571 784 605 818
rect 639 784 673 818
rect 707 784 741 818
rect 775 784 809 818
rect 843 784 877 818
rect 911 784 945 818
rect 979 784 1013 818
rect 1047 784 1081 818
rect 1115 784 1149 818
rect 1183 784 1217 818
rect 1251 784 1285 818
rect 1319 784 1353 818
rect 1387 784 1421 818
rect 1455 784 1489 818
rect 1523 784 1557 818
rect 1591 784 1625 818
rect 1659 784 1693 818
rect 1727 784 1761 818
rect 1795 784 1829 818
rect 1863 784 1897 818
rect 1931 784 1965 818
rect 1999 784 2033 818
rect 2067 784 2101 818
rect 2135 784 2169 818
rect 2203 784 2237 818
rect 2271 784 2305 818
rect 2339 784 2373 818
rect 2407 784 2441 818
rect 2475 784 2509 818
rect 2543 784 2577 818
rect 2611 784 2645 818
rect 2679 784 2713 818
rect 2747 784 2781 818
rect 2815 784 2849 818
rect 2883 784 2917 818
rect 2951 784 2985 818
rect 3019 784 3053 818
rect 3245 784 3279 818
rect 3313 784 3347 818
rect 3381 784 3415 818
rect 3449 784 3483 818
rect 3517 784 3551 818
rect 3585 784 3619 818
rect 3653 784 3687 818
rect 3721 784 3755 818
rect 3789 784 3823 818
rect 3857 784 3891 818
rect 3925 784 3959 818
rect 3993 784 4027 818
rect 4061 784 4095 818
rect 4129 784 4163 818
rect 4197 784 4231 818
rect 4265 784 4299 818
rect 4333 784 4367 818
rect 4401 784 4435 818
rect 4469 784 4503 818
rect 4537 784 4571 818
rect 4605 784 4639 818
rect 4673 784 4707 818
rect 4741 784 4775 818
rect 4809 784 4843 818
rect 4877 784 4911 818
rect 4945 784 4979 818
rect 5013 784 5047 818
rect 5081 784 5115 818
rect 5149 784 5183 818
rect 5217 784 5251 818
rect 5285 784 5319 818
rect 5353 784 5387 818
rect 5421 784 5455 818
rect 5489 784 5523 818
rect 5557 784 5591 818
rect 5625 784 5659 818
rect 5693 784 5727 818
rect 5761 784 5795 818
rect 5829 784 5863 818
rect 5897 784 5931 818
rect 5965 784 5999 818
rect 6033 784 6067 818
rect 6101 784 6135 818
rect 6169 784 6203 818
rect 9545 914 9579 948
rect 9613 914 9647 948
rect 9681 914 9715 948
rect 9749 914 9783 948
rect 9817 914 9851 948
rect 9885 914 9919 948
rect 9953 914 9987 948
rect 10021 914 10055 948
rect 10089 914 10123 948
rect 10157 914 10191 948
rect 10225 914 10259 948
rect 10293 914 10327 948
rect 10361 914 10395 948
rect 10429 914 10463 948
rect 10497 914 10531 948
rect 10565 914 10599 948
rect 10633 914 10667 948
rect 10701 914 10735 948
rect 10769 914 10803 948
rect 10837 914 10871 948
rect 10905 914 10939 948
rect 10973 914 11007 948
rect 11041 914 11075 948
rect 11109 914 11143 948
rect 11177 914 11211 948
rect 11245 914 11279 948
rect 11313 914 11347 948
rect 11381 914 11415 948
rect 11449 914 11483 948
rect 11517 914 11551 948
rect 11585 914 11619 948
rect 11653 914 11687 948
rect 11721 914 11755 948
rect 11789 914 11823 948
rect 11857 914 11891 948
rect 11925 914 11959 948
rect 11993 914 12027 948
rect 12061 914 12095 948
rect 12129 914 12163 948
rect 12197 914 12231 948
rect 12265 914 12299 948
rect 12333 914 12367 948
rect 12401 914 12435 948
rect 12469 914 12503 948
rect 12695 914 12729 948
rect 12763 914 12797 948
rect 12831 914 12865 948
rect 12899 914 12933 948
rect 12967 914 13001 948
rect 13035 914 13069 948
rect 13103 914 13137 948
rect 13171 914 13205 948
rect 13239 914 13273 948
rect 13307 914 13341 948
rect 13375 914 13409 948
rect 13443 914 13477 948
rect 13511 914 13545 948
rect 13579 914 13613 948
rect 13647 914 13681 948
rect 13715 914 13749 948
rect 13783 914 13817 948
rect 13851 914 13885 948
rect 13919 914 13953 948
rect 13987 914 14021 948
rect 14055 914 14089 948
rect 14123 914 14157 948
rect 14191 914 14225 948
rect 14259 914 14293 948
rect 14327 914 14361 948
rect 14395 914 14429 948
rect 14463 914 14497 948
rect 14531 914 14565 948
rect 14599 914 14633 948
rect 14667 914 14701 948
rect 14735 914 14769 948
rect 14803 914 14837 948
rect 14871 914 14905 948
rect 14939 914 14973 948
rect 15007 914 15041 948
rect 15075 914 15109 948
rect 15143 914 15177 948
rect 15211 914 15245 948
rect 15279 914 15313 948
rect 15347 914 15381 948
rect 15415 914 15449 948
rect 15483 914 15517 948
rect 15551 914 15585 948
rect 15619 914 15653 948
rect 15845 914 15879 948
rect 15913 914 15947 948
rect 15981 914 16015 948
rect 16049 914 16083 948
rect 16117 914 16151 948
rect 16185 914 16219 948
rect 16253 914 16287 948
rect 16321 914 16355 948
rect 16389 914 16423 948
rect 16457 914 16491 948
rect 16525 914 16559 948
rect 16593 914 16627 948
rect 16661 914 16695 948
rect 16729 914 16763 948
rect 16797 914 16831 948
rect 16865 914 16899 948
rect 16933 914 16967 948
rect 17001 914 17035 948
rect 17069 914 17103 948
rect 17137 914 17171 948
rect 17205 914 17239 948
rect 17273 914 17307 948
rect 17341 914 17375 948
rect 17409 914 17443 948
rect 17477 914 17511 948
rect 17545 914 17579 948
rect 17613 914 17647 948
rect 17681 914 17715 948
rect 17749 914 17783 948
rect 17817 914 17851 948
rect 17885 914 17919 948
rect 17953 914 17987 948
rect 18021 914 18055 948
rect 18089 914 18123 948
rect 18157 914 18191 948
rect 18225 914 18259 948
rect 18293 914 18327 948
rect 18361 914 18395 948
rect 18429 914 18463 948
rect 18497 914 18531 948
rect 18565 914 18599 948
rect 18633 914 18667 948
rect 18701 914 18735 948
rect 18769 914 18803 948
rect 18995 914 19029 948
rect 19063 914 19097 948
rect 19131 914 19165 948
rect 19199 914 19233 948
rect 19267 914 19301 948
rect 19335 914 19369 948
rect 19403 914 19437 948
rect 19471 914 19505 948
rect 19539 914 19573 948
rect 19607 914 19641 948
rect 19675 914 19709 948
rect 19743 914 19777 948
rect 19811 914 19845 948
rect 19879 914 19913 948
rect 19947 914 19981 948
rect 20015 914 20049 948
rect 20083 914 20117 948
rect 20151 914 20185 948
rect 20219 914 20253 948
rect 20287 914 20321 948
rect 20355 914 20389 948
rect 20423 914 20457 948
rect 20491 914 20525 948
rect 20559 914 20593 948
rect 20627 914 20661 948
rect 20695 914 20729 948
rect 20763 914 20797 948
rect 20831 914 20865 948
rect 20899 914 20933 948
rect 20967 914 21001 948
rect 21035 914 21069 948
rect 21103 914 21137 948
rect 21171 914 21205 948
rect 21239 914 21273 948
rect 21307 914 21341 948
rect 21375 914 21409 948
rect 21443 914 21477 948
rect 21511 914 21545 948
rect 21579 914 21613 948
rect 21647 914 21681 948
rect 21715 914 21749 948
rect 21783 914 21817 948
rect 21851 914 21885 948
rect 21919 914 21953 948
rect 6395 758 6429 792
rect 6463 758 6497 792
rect 6531 758 6565 792
rect 6599 758 6633 792
rect 6667 758 6701 792
rect 6735 758 6769 792
rect 6803 758 6837 792
rect 6871 758 6905 792
rect 6939 758 6973 792
rect 7007 758 7041 792
rect 7075 758 7109 792
rect 7143 758 7177 792
rect 7211 758 7245 792
rect 7279 758 7313 792
rect 7347 758 7381 792
rect 7415 758 7449 792
rect 7483 758 7517 792
rect 7551 758 7585 792
rect 7619 758 7653 792
rect 7687 758 7721 792
rect 7755 758 7789 792
rect 7823 758 7857 792
rect 7891 758 7925 792
rect 7959 758 7993 792
rect 8027 758 8061 792
rect 8095 758 8129 792
rect 8163 758 8197 792
rect 8231 758 8265 792
rect 8299 758 8333 792
rect 8367 758 8401 792
rect 8435 758 8469 792
rect 8503 758 8537 792
rect 8571 758 8605 792
rect 8639 758 8673 792
rect 8707 758 8741 792
rect 8775 758 8809 792
rect 8843 758 8877 792
rect 8911 758 8945 792
rect 8979 758 9013 792
rect 9047 758 9081 792
rect 9115 758 9149 792
rect 9183 758 9217 792
rect 9251 758 9285 792
rect 9319 758 9353 792
rect 95 628 129 662
rect 163 628 197 662
rect 231 628 265 662
rect 299 628 333 662
rect 367 628 401 662
rect 435 628 469 662
rect 503 628 537 662
rect 571 628 605 662
rect 639 628 673 662
rect 707 628 741 662
rect 775 628 809 662
rect 843 628 877 662
rect 911 628 945 662
rect 979 628 1013 662
rect 1047 628 1081 662
rect 1115 628 1149 662
rect 1183 628 1217 662
rect 1251 628 1285 662
rect 1319 628 1353 662
rect 1387 628 1421 662
rect 1455 628 1489 662
rect 1523 628 1557 662
rect 1591 628 1625 662
rect 1659 628 1693 662
rect 1727 628 1761 662
rect 1795 628 1829 662
rect 1863 628 1897 662
rect 1931 628 1965 662
rect 1999 628 2033 662
rect 2067 628 2101 662
rect 2135 628 2169 662
rect 2203 628 2237 662
rect 2271 628 2305 662
rect 2339 628 2373 662
rect 2407 628 2441 662
rect 2475 628 2509 662
rect 2543 628 2577 662
rect 2611 628 2645 662
rect 2679 628 2713 662
rect 2747 628 2781 662
rect 2815 628 2849 662
rect 2883 628 2917 662
rect 2951 628 2985 662
rect 3019 628 3053 662
rect 3245 628 3279 662
rect 3313 628 3347 662
rect 3381 628 3415 662
rect 3449 628 3483 662
rect 3517 628 3551 662
rect 3585 628 3619 662
rect 3653 628 3687 662
rect 3721 628 3755 662
rect 3789 628 3823 662
rect 3857 628 3891 662
rect 3925 628 3959 662
rect 3993 628 4027 662
rect 4061 628 4095 662
rect 4129 628 4163 662
rect 4197 628 4231 662
rect 4265 628 4299 662
rect 4333 628 4367 662
rect 4401 628 4435 662
rect 4469 628 4503 662
rect 4537 628 4571 662
rect 4605 628 4639 662
rect 4673 628 4707 662
rect 4741 628 4775 662
rect 4809 628 4843 662
rect 4877 628 4911 662
rect 4945 628 4979 662
rect 5013 628 5047 662
rect 5081 628 5115 662
rect 5149 628 5183 662
rect 5217 628 5251 662
rect 5285 628 5319 662
rect 5353 628 5387 662
rect 5421 628 5455 662
rect 5489 628 5523 662
rect 5557 628 5591 662
rect 5625 628 5659 662
rect 5693 628 5727 662
rect 5761 628 5795 662
rect 5829 628 5863 662
rect 5897 628 5931 662
rect 5965 628 5999 662
rect 6033 628 6067 662
rect 6101 628 6135 662
rect 6169 628 6203 662
rect 9545 758 9579 792
rect 9613 758 9647 792
rect 9681 758 9715 792
rect 9749 758 9783 792
rect 9817 758 9851 792
rect 9885 758 9919 792
rect 9953 758 9987 792
rect 10021 758 10055 792
rect 10089 758 10123 792
rect 10157 758 10191 792
rect 10225 758 10259 792
rect 10293 758 10327 792
rect 10361 758 10395 792
rect 10429 758 10463 792
rect 10497 758 10531 792
rect 10565 758 10599 792
rect 10633 758 10667 792
rect 10701 758 10735 792
rect 10769 758 10803 792
rect 10837 758 10871 792
rect 10905 758 10939 792
rect 10973 758 11007 792
rect 11041 758 11075 792
rect 11109 758 11143 792
rect 11177 758 11211 792
rect 11245 758 11279 792
rect 11313 758 11347 792
rect 11381 758 11415 792
rect 11449 758 11483 792
rect 11517 758 11551 792
rect 11585 758 11619 792
rect 11653 758 11687 792
rect 11721 758 11755 792
rect 11789 758 11823 792
rect 11857 758 11891 792
rect 11925 758 11959 792
rect 11993 758 12027 792
rect 12061 758 12095 792
rect 12129 758 12163 792
rect 12197 758 12231 792
rect 12265 758 12299 792
rect 12333 758 12367 792
rect 12401 758 12435 792
rect 12469 758 12503 792
rect 12695 758 12729 792
rect 12763 758 12797 792
rect 12831 758 12865 792
rect 12899 758 12933 792
rect 12967 758 13001 792
rect 13035 758 13069 792
rect 13103 758 13137 792
rect 13171 758 13205 792
rect 13239 758 13273 792
rect 13307 758 13341 792
rect 13375 758 13409 792
rect 13443 758 13477 792
rect 13511 758 13545 792
rect 13579 758 13613 792
rect 13647 758 13681 792
rect 13715 758 13749 792
rect 13783 758 13817 792
rect 13851 758 13885 792
rect 13919 758 13953 792
rect 13987 758 14021 792
rect 14055 758 14089 792
rect 14123 758 14157 792
rect 14191 758 14225 792
rect 14259 758 14293 792
rect 14327 758 14361 792
rect 14395 758 14429 792
rect 14463 758 14497 792
rect 14531 758 14565 792
rect 14599 758 14633 792
rect 14667 758 14701 792
rect 14735 758 14769 792
rect 14803 758 14837 792
rect 14871 758 14905 792
rect 14939 758 14973 792
rect 15007 758 15041 792
rect 15075 758 15109 792
rect 15143 758 15177 792
rect 15211 758 15245 792
rect 15279 758 15313 792
rect 15347 758 15381 792
rect 15415 758 15449 792
rect 15483 758 15517 792
rect 15551 758 15585 792
rect 15619 758 15653 792
rect 15845 758 15879 792
rect 15913 758 15947 792
rect 15981 758 16015 792
rect 16049 758 16083 792
rect 16117 758 16151 792
rect 16185 758 16219 792
rect 16253 758 16287 792
rect 16321 758 16355 792
rect 16389 758 16423 792
rect 16457 758 16491 792
rect 16525 758 16559 792
rect 16593 758 16627 792
rect 16661 758 16695 792
rect 16729 758 16763 792
rect 16797 758 16831 792
rect 16865 758 16899 792
rect 16933 758 16967 792
rect 17001 758 17035 792
rect 17069 758 17103 792
rect 17137 758 17171 792
rect 17205 758 17239 792
rect 17273 758 17307 792
rect 17341 758 17375 792
rect 17409 758 17443 792
rect 17477 758 17511 792
rect 17545 758 17579 792
rect 17613 758 17647 792
rect 17681 758 17715 792
rect 17749 758 17783 792
rect 17817 758 17851 792
rect 17885 758 17919 792
rect 17953 758 17987 792
rect 18021 758 18055 792
rect 18089 758 18123 792
rect 18157 758 18191 792
rect 18225 758 18259 792
rect 18293 758 18327 792
rect 18361 758 18395 792
rect 18429 758 18463 792
rect 18497 758 18531 792
rect 18565 758 18599 792
rect 18633 758 18667 792
rect 18701 758 18735 792
rect 18769 758 18803 792
rect 18995 758 19029 792
rect 19063 758 19097 792
rect 19131 758 19165 792
rect 19199 758 19233 792
rect 19267 758 19301 792
rect 19335 758 19369 792
rect 19403 758 19437 792
rect 19471 758 19505 792
rect 19539 758 19573 792
rect 19607 758 19641 792
rect 19675 758 19709 792
rect 19743 758 19777 792
rect 19811 758 19845 792
rect 19879 758 19913 792
rect 19947 758 19981 792
rect 20015 758 20049 792
rect 20083 758 20117 792
rect 20151 758 20185 792
rect 20219 758 20253 792
rect 20287 758 20321 792
rect 20355 758 20389 792
rect 20423 758 20457 792
rect 20491 758 20525 792
rect 20559 758 20593 792
rect 20627 758 20661 792
rect 20695 758 20729 792
rect 20763 758 20797 792
rect 20831 758 20865 792
rect 20899 758 20933 792
rect 20967 758 21001 792
rect 21035 758 21069 792
rect 21103 758 21137 792
rect 21171 758 21205 792
rect 21239 758 21273 792
rect 21307 758 21341 792
rect 21375 758 21409 792
rect 21443 758 21477 792
rect 21511 758 21545 792
rect 21579 758 21613 792
rect 21647 758 21681 792
rect 21715 758 21749 792
rect 21783 758 21817 792
rect 21851 758 21885 792
rect 21919 758 21953 792
rect 22390 1136 22424 1170
rect 22458 1136 22492 1170
rect 22526 1136 22560 1170
rect 22594 1136 22628 1170
rect 22662 1136 22696 1170
rect 22730 1136 22764 1170
rect 22798 1136 22832 1170
rect 22866 1136 22900 1170
rect 22934 1136 22968 1170
rect 23002 1136 23036 1170
rect 23070 1136 23104 1170
rect 23138 1136 23172 1170
rect 23206 1136 23240 1170
rect 23274 1136 23308 1170
rect 23342 1136 23376 1170
rect 23410 1136 23444 1170
rect 23478 1136 23512 1170
rect 23546 1136 23580 1170
rect 23614 1136 23648 1170
rect 23682 1136 23716 1170
rect 23750 1136 23784 1170
rect 23818 1136 23852 1170
rect 23886 1136 23920 1170
rect 23954 1136 23988 1170
rect 24022 1136 24056 1170
rect 24090 1136 24124 1170
rect 24158 1136 24192 1170
rect 24226 1136 24260 1170
rect 24294 1136 24328 1170
rect 22390 980 22424 1014
rect 22458 980 22492 1014
rect 22526 980 22560 1014
rect 22594 980 22628 1014
rect 22662 980 22696 1014
rect 22730 980 22764 1014
rect 22798 980 22832 1014
rect 22866 980 22900 1014
rect 22934 980 22968 1014
rect 23002 980 23036 1014
rect 23070 980 23104 1014
rect 23138 980 23172 1014
rect 23206 980 23240 1014
rect 23274 980 23308 1014
rect 23342 980 23376 1014
rect 23410 980 23444 1014
rect 23478 980 23512 1014
rect 23546 980 23580 1014
rect 23614 980 23648 1014
rect 23682 980 23716 1014
rect 23750 980 23784 1014
rect 23818 980 23852 1014
rect 23886 980 23920 1014
rect 23954 980 23988 1014
rect 24022 980 24056 1014
rect 24090 980 24124 1014
rect 24158 980 24192 1014
rect 24226 980 24260 1014
rect 24294 980 24328 1014
rect 22390 824 22424 858
rect 22458 824 22492 858
rect 22526 824 22560 858
rect 22594 824 22628 858
rect 22662 824 22696 858
rect 22730 824 22764 858
rect 22798 824 22832 858
rect 22866 824 22900 858
rect 22934 824 22968 858
rect 23002 824 23036 858
rect 23070 824 23104 858
rect 23138 824 23172 858
rect 23206 824 23240 858
rect 23274 824 23308 858
rect 23342 824 23376 858
rect 23410 824 23444 858
rect 23478 824 23512 858
rect 23546 824 23580 858
rect 23614 824 23648 858
rect 23682 824 23716 858
rect 23750 824 23784 858
rect 23818 824 23852 858
rect 23886 824 23920 858
rect 23954 824 23988 858
rect 24022 824 24056 858
rect 24090 824 24124 858
rect 24158 824 24192 858
rect 24226 824 24260 858
rect 24294 824 24328 858
rect 22390 668 22424 702
rect 22458 668 22492 702
rect 22526 668 22560 702
rect 22594 668 22628 702
rect 22662 668 22696 702
rect 22730 668 22764 702
rect 22798 668 22832 702
rect 22866 668 22900 702
rect 22934 668 22968 702
rect 23002 668 23036 702
rect 23070 668 23104 702
rect 23138 668 23172 702
rect 23206 668 23240 702
rect 23274 668 23308 702
rect 23342 668 23376 702
rect 23410 668 23444 702
rect 23478 668 23512 702
rect 23546 668 23580 702
rect 23614 668 23648 702
rect 23682 668 23716 702
rect 23750 668 23784 702
rect 23818 668 23852 702
rect 23886 668 23920 702
rect 23954 668 23988 702
rect 24022 668 24056 702
rect 24090 668 24124 702
rect 24158 668 24192 702
rect 24226 668 24260 702
rect 24294 668 24328 702
rect 6395 602 6429 636
rect 6463 602 6497 636
rect 6531 602 6565 636
rect 6599 602 6633 636
rect 6667 602 6701 636
rect 6735 602 6769 636
rect 6803 602 6837 636
rect 6871 602 6905 636
rect 6939 602 6973 636
rect 7007 602 7041 636
rect 7075 602 7109 636
rect 7143 602 7177 636
rect 7211 602 7245 636
rect 7279 602 7313 636
rect 7347 602 7381 636
rect 7415 602 7449 636
rect 7483 602 7517 636
rect 7551 602 7585 636
rect 7619 602 7653 636
rect 7687 602 7721 636
rect 7755 602 7789 636
rect 7823 602 7857 636
rect 7891 602 7925 636
rect 7959 602 7993 636
rect 8027 602 8061 636
rect 8095 602 8129 636
rect 8163 602 8197 636
rect 8231 602 8265 636
rect 8299 602 8333 636
rect 8367 602 8401 636
rect 8435 602 8469 636
rect 8503 602 8537 636
rect 8571 602 8605 636
rect 8639 602 8673 636
rect 8707 602 8741 636
rect 8775 602 8809 636
rect 8843 602 8877 636
rect 8911 602 8945 636
rect 8979 602 9013 636
rect 9047 602 9081 636
rect 9115 602 9149 636
rect 9183 602 9217 636
rect 9251 602 9285 636
rect 9319 602 9353 636
rect 9545 602 9579 636
rect 9613 602 9647 636
rect 9681 602 9715 636
rect 9749 602 9783 636
rect 9817 602 9851 636
rect 9885 602 9919 636
rect 9953 602 9987 636
rect 10021 602 10055 636
rect 10089 602 10123 636
rect 10157 602 10191 636
rect 10225 602 10259 636
rect 10293 602 10327 636
rect 10361 602 10395 636
rect 10429 602 10463 636
rect 10497 602 10531 636
rect 10565 602 10599 636
rect 10633 602 10667 636
rect 10701 602 10735 636
rect 10769 602 10803 636
rect 10837 602 10871 636
rect 10905 602 10939 636
rect 10973 602 11007 636
rect 11041 602 11075 636
rect 11109 602 11143 636
rect 11177 602 11211 636
rect 11245 602 11279 636
rect 11313 602 11347 636
rect 11381 602 11415 636
rect 11449 602 11483 636
rect 11517 602 11551 636
rect 11585 602 11619 636
rect 11653 602 11687 636
rect 11721 602 11755 636
rect 11789 602 11823 636
rect 11857 602 11891 636
rect 11925 602 11959 636
rect 11993 602 12027 636
rect 12061 602 12095 636
rect 12129 602 12163 636
rect 12197 602 12231 636
rect 12265 602 12299 636
rect 12333 602 12367 636
rect 12401 602 12435 636
rect 12469 602 12503 636
rect 12695 602 12729 636
rect 12763 602 12797 636
rect 12831 602 12865 636
rect 12899 602 12933 636
rect 12967 602 13001 636
rect 13035 602 13069 636
rect 13103 602 13137 636
rect 13171 602 13205 636
rect 13239 602 13273 636
rect 13307 602 13341 636
rect 13375 602 13409 636
rect 13443 602 13477 636
rect 13511 602 13545 636
rect 13579 602 13613 636
rect 13647 602 13681 636
rect 13715 602 13749 636
rect 13783 602 13817 636
rect 13851 602 13885 636
rect 13919 602 13953 636
rect 13987 602 14021 636
rect 14055 602 14089 636
rect 14123 602 14157 636
rect 14191 602 14225 636
rect 14259 602 14293 636
rect 14327 602 14361 636
rect 14395 602 14429 636
rect 14463 602 14497 636
rect 14531 602 14565 636
rect 14599 602 14633 636
rect 14667 602 14701 636
rect 14735 602 14769 636
rect 14803 602 14837 636
rect 14871 602 14905 636
rect 14939 602 14973 636
rect 15007 602 15041 636
rect 15075 602 15109 636
rect 15143 602 15177 636
rect 15211 602 15245 636
rect 15279 602 15313 636
rect 15347 602 15381 636
rect 15415 602 15449 636
rect 15483 602 15517 636
rect 15551 602 15585 636
rect 15619 602 15653 636
rect 15845 602 15879 636
rect 15913 602 15947 636
rect 15981 602 16015 636
rect 16049 602 16083 636
rect 16117 602 16151 636
rect 16185 602 16219 636
rect 16253 602 16287 636
rect 16321 602 16355 636
rect 16389 602 16423 636
rect 16457 602 16491 636
rect 16525 602 16559 636
rect 16593 602 16627 636
rect 16661 602 16695 636
rect 16729 602 16763 636
rect 16797 602 16831 636
rect 16865 602 16899 636
rect 16933 602 16967 636
rect 17001 602 17035 636
rect 17069 602 17103 636
rect 17137 602 17171 636
rect 17205 602 17239 636
rect 17273 602 17307 636
rect 17341 602 17375 636
rect 17409 602 17443 636
rect 17477 602 17511 636
rect 17545 602 17579 636
rect 17613 602 17647 636
rect 17681 602 17715 636
rect 17749 602 17783 636
rect 17817 602 17851 636
rect 17885 602 17919 636
rect 17953 602 17987 636
rect 18021 602 18055 636
rect 18089 602 18123 636
rect 18157 602 18191 636
rect 18225 602 18259 636
rect 18293 602 18327 636
rect 18361 602 18395 636
rect 18429 602 18463 636
rect 18497 602 18531 636
rect 18565 602 18599 636
rect 18633 602 18667 636
rect 18701 602 18735 636
rect 18769 602 18803 636
rect 18995 602 19029 636
rect 19063 602 19097 636
rect 19131 602 19165 636
rect 19199 602 19233 636
rect 19267 602 19301 636
rect 19335 602 19369 636
rect 19403 602 19437 636
rect 19471 602 19505 636
rect 19539 602 19573 636
rect 19607 602 19641 636
rect 19675 602 19709 636
rect 19743 602 19777 636
rect 19811 602 19845 636
rect 19879 602 19913 636
rect 19947 602 19981 636
rect 20015 602 20049 636
rect 20083 602 20117 636
rect 20151 602 20185 636
rect 20219 602 20253 636
rect 20287 602 20321 636
rect 20355 602 20389 636
rect 20423 602 20457 636
rect 20491 602 20525 636
rect 20559 602 20593 636
rect 20627 602 20661 636
rect 20695 602 20729 636
rect 20763 602 20797 636
rect 20831 602 20865 636
rect 20899 602 20933 636
rect 20967 602 21001 636
rect 21035 602 21069 636
rect 21103 602 21137 636
rect 21171 602 21205 636
rect 21239 602 21273 636
rect 21307 602 21341 636
rect 21375 602 21409 636
rect 21443 602 21477 636
rect 21511 602 21545 636
rect 21579 602 21613 636
rect 21647 602 21681 636
rect 21715 602 21749 636
rect 21783 602 21817 636
rect 21851 602 21885 636
rect 21919 602 21953 636
<< poly >>
rect 22216 2045 22340 2061
rect 22216 2011 22248 2045
rect 22282 2011 22340 2045
rect 22216 1974 22340 2011
rect 22216 1940 22248 1974
rect 22282 1961 22340 1974
rect 24340 1961 24366 2061
rect 22282 1940 22314 1961
rect 22216 1905 22314 1940
rect 22216 1903 22340 1905
rect 22216 1869 22248 1903
rect 22282 1869 22340 1903
rect 22216 1832 22340 1869
rect 22216 1798 22248 1832
rect 22282 1805 22340 1832
rect 24340 1805 24366 1905
rect 22282 1798 22314 1805
rect 22216 1761 22314 1798
rect 22216 1727 22248 1761
rect 22282 1749 22314 1761
rect 22282 1727 22340 1749
rect 22216 1690 22340 1727
rect 22216 1656 22248 1690
rect 22282 1656 22340 1690
rect 22216 1649 22340 1656
rect 24340 1649 24366 1749
rect 22216 1619 22314 1649
rect 22216 1585 22248 1619
rect 22282 1593 22314 1619
rect 22282 1585 22340 1593
rect 22216 1548 22340 1585
rect 22216 1514 22248 1548
rect 22282 1514 22340 1548
rect 22216 1493 22340 1514
rect 24340 1493 24366 1593
rect 22216 1477 22314 1493
rect 22216 1443 22248 1477
rect 22282 1443 22314 1477
rect 22216 1437 22314 1443
rect 22216 1406 22340 1437
rect 22216 1372 22248 1406
rect 22282 1372 22340 1406
rect 22216 1337 22340 1372
rect 24340 1337 24366 1437
rect 22216 1335 22314 1337
rect 22216 1301 22248 1335
rect 22282 1301 22314 1335
rect 22216 1281 22314 1301
rect 22216 1264 22340 1281
rect 22216 1230 22248 1264
rect 22282 1230 22340 1264
rect 6241 1193 6365 1215
rect 6241 1159 6273 1193
rect 6307 1159 6365 1193
rect 6241 1115 6365 1159
rect 9365 1199 9515 1215
rect 9365 1165 9423 1199
rect 9457 1165 9515 1199
rect 9365 1128 9515 1165
rect 9365 1115 9423 1128
rect 6241 1081 6273 1115
rect 6307 1081 6339 1115
rect 6241 1059 6339 1081
rect 9391 1094 9423 1115
rect 9457 1115 9515 1128
rect 12515 1199 12665 1215
rect 12515 1165 12573 1199
rect 12607 1165 12665 1199
rect 12515 1128 12665 1165
rect 12515 1115 12573 1128
rect 9457 1094 9489 1115
rect 9391 1059 9489 1094
rect 12541 1094 12573 1115
rect 12607 1115 12665 1128
rect 15665 1199 15815 1215
rect 15665 1165 15723 1199
rect 15757 1165 15815 1199
rect 15665 1128 15815 1165
rect 15665 1115 15723 1128
rect 12607 1094 12639 1115
rect 12541 1059 12639 1094
rect 15691 1094 15723 1115
rect 15757 1115 15815 1128
rect 18815 1199 18965 1215
rect 18815 1165 18873 1199
rect 18907 1165 18965 1199
rect 18815 1128 18965 1165
rect 18815 1115 18873 1128
rect 15757 1094 15789 1115
rect 15691 1059 15789 1094
rect 18841 1094 18873 1115
rect 18907 1115 18965 1128
rect 21965 1199 22089 1215
rect 21965 1165 22023 1199
rect 22057 1165 22089 1199
rect 21965 1128 22089 1165
rect 21965 1115 22023 1128
rect 18907 1094 18939 1115
rect 18841 1059 18939 1094
rect 21991 1094 22023 1115
rect 22057 1094 22089 1128
rect 21991 1059 22089 1094
rect 6241 1037 6365 1059
rect 6241 1003 6273 1037
rect 6307 1003 6365 1037
rect 6241 959 6365 1003
rect 9365 1057 9515 1059
rect 9365 1023 9423 1057
rect 9457 1023 9515 1057
rect 9365 985 9515 1023
rect 9365 959 9423 985
rect 6241 925 6273 959
rect 6307 925 6339 959
rect 6241 903 6339 925
rect 9391 951 9423 959
rect 9457 959 9515 985
rect 12515 1057 12665 1059
rect 12515 1023 12573 1057
rect 12607 1023 12665 1057
rect 12515 985 12665 1023
rect 12515 959 12573 985
rect 9457 951 9489 959
rect 9391 913 9489 951
rect 9391 903 9423 913
rect 6241 881 6365 903
rect 6241 847 6273 881
rect 6307 847 6365 881
rect 3107 794 3173 810
rect 3107 773 3123 794
rect 39 673 65 773
rect 3065 760 3123 773
rect 3157 773 3173 794
rect 6241 803 6365 847
rect 9365 879 9423 903
rect 9457 903 9489 913
rect 12541 951 12573 959
rect 12607 959 12665 985
rect 15665 1057 15815 1059
rect 15665 1023 15723 1057
rect 15757 1023 15815 1057
rect 15665 985 15815 1023
rect 15665 959 15723 985
rect 12607 951 12639 959
rect 12541 913 12639 951
rect 12541 903 12573 913
rect 9457 879 9515 903
rect 9365 841 9515 879
rect 9365 807 9423 841
rect 9457 807 9515 841
rect 9365 803 9515 807
rect 12515 879 12573 903
rect 12607 903 12639 913
rect 15691 951 15723 959
rect 15757 959 15815 985
rect 18815 1057 18965 1059
rect 18815 1023 18873 1057
rect 18907 1023 18965 1057
rect 18815 985 18965 1023
rect 18815 959 18873 985
rect 15757 951 15789 959
rect 15691 913 15789 951
rect 15691 903 15723 913
rect 12607 879 12665 903
rect 12515 841 12665 879
rect 12515 807 12573 841
rect 12607 807 12665 841
rect 12515 803 12665 807
rect 15665 879 15723 903
rect 15757 903 15789 913
rect 18841 951 18873 959
rect 18907 959 18965 985
rect 21965 1057 22089 1059
rect 21965 1023 22023 1057
rect 22057 1023 22089 1057
rect 21965 985 22089 1023
rect 21965 959 22023 985
rect 18907 951 18939 959
rect 18841 913 18939 951
rect 18841 903 18873 913
rect 15757 879 15815 903
rect 15665 841 15815 879
rect 15665 807 15723 841
rect 15757 807 15815 841
rect 15665 803 15815 807
rect 18815 879 18873 903
rect 18907 903 18939 913
rect 21991 951 22023 959
rect 22057 951 22089 985
rect 21991 913 22089 951
rect 21991 903 22023 913
rect 18907 879 18965 903
rect 18815 841 18965 879
rect 18815 807 18873 841
rect 18907 807 18965 841
rect 18815 803 18965 807
rect 21965 879 22023 903
rect 22057 879 22089 913
rect 21965 841 22089 879
rect 21965 807 22023 841
rect 22057 807 22089 841
rect 21965 803 22089 807
rect 6241 802 6339 803
rect 6241 773 6273 802
rect 3157 760 3215 773
rect 3065 723 3215 760
rect 3065 689 3123 723
rect 3157 689 3215 723
rect 3065 673 3215 689
rect 6215 768 6273 773
rect 6307 768 6339 802
rect 6215 747 6339 768
rect 9391 769 9489 803
rect 9391 747 9423 769
rect 6215 723 6365 747
rect 6215 689 6273 723
rect 6307 689 6365 723
rect 6215 673 6365 689
rect 6241 647 6365 673
rect 9365 735 9423 747
rect 9457 747 9489 769
rect 12541 769 12639 803
rect 12541 747 12573 769
rect 9457 735 9515 747
rect 9365 697 9515 735
rect 9365 663 9423 697
rect 9457 663 9515 697
rect 9365 647 9515 663
rect 12515 735 12573 747
rect 12607 747 12639 769
rect 15691 769 15789 803
rect 15691 747 15723 769
rect 12607 735 12665 747
rect 12515 697 12665 735
rect 12515 663 12573 697
rect 12607 663 12665 697
rect 12515 647 12665 663
rect 15665 735 15723 747
rect 15757 747 15789 769
rect 18841 769 18939 803
rect 18841 747 18873 769
rect 15757 735 15815 747
rect 15665 697 15815 735
rect 15665 663 15723 697
rect 15757 663 15815 697
rect 15665 647 15815 663
rect 18815 735 18873 747
rect 18907 747 18939 769
rect 21991 769 22089 803
rect 21991 747 22023 769
rect 18907 735 18965 747
rect 18815 697 18965 735
rect 18815 663 18873 697
rect 18907 663 18965 697
rect 18815 647 18965 663
rect 21965 735 22023 747
rect 22057 735 22089 769
rect 21965 697 22089 735
rect 22216 1193 22340 1230
rect 22216 1159 22248 1193
rect 22282 1181 22340 1193
rect 24340 1181 24366 1281
rect 22282 1159 22314 1181
rect 22216 1125 22314 1159
rect 22216 1122 22340 1125
rect 22216 1088 22248 1122
rect 22282 1088 22340 1122
rect 22216 1051 22340 1088
rect 22216 1017 22248 1051
rect 22282 1025 22340 1051
rect 24340 1025 24366 1125
rect 22282 1017 22314 1025
rect 22216 979 22314 1017
rect 22216 945 22248 979
rect 22282 969 22314 979
rect 22282 945 22340 969
rect 22216 907 22340 945
rect 22216 873 22248 907
rect 22282 873 22340 907
rect 22216 869 22340 873
rect 24340 869 24366 969
rect 22216 835 22314 869
rect 22216 801 22248 835
rect 22282 813 22314 835
rect 22282 801 22340 813
rect 22216 763 22340 801
rect 22216 729 22248 763
rect 22282 729 22340 763
rect 22216 713 22340 729
rect 24340 713 24366 813
rect 21965 663 22023 697
rect 22057 663 22089 697
rect 21965 647 22089 663
<< polycont >>
rect 22248 2011 22282 2045
rect 22248 1940 22282 1974
rect 22248 1869 22282 1903
rect 22248 1798 22282 1832
rect 22248 1727 22282 1761
rect 22248 1656 22282 1690
rect 22248 1585 22282 1619
rect 22248 1514 22282 1548
rect 22248 1443 22282 1477
rect 22248 1372 22282 1406
rect 22248 1301 22282 1335
rect 22248 1230 22282 1264
rect 6273 1159 6307 1193
rect 9423 1165 9457 1199
rect 6273 1081 6307 1115
rect 9423 1094 9457 1128
rect 12573 1165 12607 1199
rect 12573 1094 12607 1128
rect 15723 1165 15757 1199
rect 15723 1094 15757 1128
rect 18873 1165 18907 1199
rect 18873 1094 18907 1128
rect 22023 1165 22057 1199
rect 22023 1094 22057 1128
rect 6273 1003 6307 1037
rect 9423 1023 9457 1057
rect 6273 925 6307 959
rect 9423 951 9457 985
rect 12573 1023 12607 1057
rect 6273 847 6307 881
rect 3123 760 3157 794
rect 9423 879 9457 913
rect 12573 951 12607 985
rect 15723 1023 15757 1057
rect 9423 807 9457 841
rect 12573 879 12607 913
rect 15723 951 15757 985
rect 18873 1023 18907 1057
rect 12573 807 12607 841
rect 15723 879 15757 913
rect 18873 951 18907 985
rect 22023 1023 22057 1057
rect 15723 807 15757 841
rect 18873 879 18907 913
rect 22023 951 22057 985
rect 18873 807 18907 841
rect 22023 879 22057 913
rect 22023 807 22057 841
rect 3123 689 3157 723
rect 6273 768 6307 802
rect 6273 689 6307 723
rect 9423 735 9457 769
rect 9423 663 9457 697
rect 12573 735 12607 769
rect 12573 663 12607 697
rect 15723 735 15757 769
rect 15723 663 15757 697
rect 18873 735 18907 769
rect 18873 663 18907 697
rect 22023 735 22057 769
rect 22248 1159 22282 1193
rect 22248 1088 22282 1122
rect 22248 1017 22282 1051
rect 22248 945 22282 979
rect 22248 873 22282 907
rect 22248 801 22282 835
rect 22248 729 22282 763
rect 22023 663 22057 697
<< locali >>
rect 22424 2072 22438 2106
rect 22492 2072 22510 2106
rect 22560 2072 22582 2106
rect 22628 2072 22654 2106
rect 22696 2072 22726 2106
rect 22764 2072 22798 2106
rect 22832 2072 22866 2106
rect 22904 2072 22934 2106
rect 22976 2072 23002 2106
rect 23048 2072 23070 2106
rect 23120 2072 23138 2106
rect 23192 2072 23206 2106
rect 23264 2072 23274 2106
rect 23336 2072 23342 2106
rect 23408 2072 23410 2106
rect 23444 2072 23446 2106
rect 23512 2072 23518 2106
rect 23580 2072 23590 2106
rect 23648 2072 23662 2106
rect 23716 2072 23734 2106
rect 23784 2072 23806 2106
rect 23852 2072 23878 2106
rect 23920 2072 23950 2106
rect 23988 2072 24022 2106
rect 24056 2072 24090 2106
rect 24128 2072 24158 2106
rect 24200 2072 24226 2106
rect 24272 2072 24294 2106
rect 22248 2049 22282 2061
rect 22248 1974 22282 2011
rect 22248 1903 22282 1940
rect 22424 1916 22438 1950
rect 22492 1916 22510 1950
rect 22560 1916 22582 1950
rect 22628 1916 22654 1950
rect 22696 1916 22726 1950
rect 22764 1916 22798 1950
rect 22832 1916 22866 1950
rect 22904 1916 22934 1950
rect 22976 1916 23002 1950
rect 23048 1916 23070 1950
rect 23120 1916 23138 1950
rect 23192 1916 23206 1950
rect 23264 1916 23274 1950
rect 23336 1916 23342 1950
rect 23408 1916 23410 1950
rect 23444 1916 23446 1950
rect 23512 1916 23518 1950
rect 23580 1916 23590 1950
rect 23648 1916 23662 1950
rect 23716 1916 23734 1950
rect 23784 1916 23806 1950
rect 23852 1916 23878 1950
rect 23920 1916 23950 1950
rect 23988 1916 24022 1950
rect 24056 1916 24090 1950
rect 24128 1916 24158 1950
rect 24200 1916 24226 1950
rect 24272 1916 24294 1950
rect 22248 1832 22282 1865
rect 22248 1761 22282 1790
rect 22424 1760 22438 1794
rect 22492 1760 22510 1794
rect 22560 1760 22582 1794
rect 22628 1760 22654 1794
rect 22696 1760 22726 1794
rect 22764 1760 22798 1794
rect 22832 1760 22866 1794
rect 22904 1760 22934 1794
rect 22976 1760 23002 1794
rect 23048 1760 23070 1794
rect 23120 1760 23138 1794
rect 23192 1760 23206 1794
rect 23264 1760 23274 1794
rect 23336 1760 23342 1794
rect 23408 1760 23410 1794
rect 23444 1760 23446 1794
rect 23512 1760 23518 1794
rect 23580 1760 23590 1794
rect 23648 1760 23662 1794
rect 23716 1760 23734 1794
rect 23784 1760 23806 1794
rect 23852 1760 23878 1794
rect 23920 1760 23950 1794
rect 23988 1760 24022 1794
rect 24056 1760 24090 1794
rect 24128 1760 24158 1794
rect 24200 1760 24226 1794
rect 24272 1760 24294 1794
rect 22248 1690 22282 1714
rect 22248 1619 22282 1638
rect 22424 1604 22438 1638
rect 22492 1604 22510 1638
rect 22560 1604 22582 1638
rect 22628 1604 22654 1638
rect 22696 1604 22726 1638
rect 22764 1604 22798 1638
rect 22832 1604 22866 1638
rect 22904 1604 22934 1638
rect 22976 1604 23002 1638
rect 23048 1604 23070 1638
rect 23120 1604 23138 1638
rect 23192 1604 23206 1638
rect 23264 1604 23274 1638
rect 23336 1604 23342 1638
rect 23408 1604 23410 1638
rect 23444 1604 23446 1638
rect 23512 1604 23518 1638
rect 23580 1604 23590 1638
rect 23648 1604 23662 1638
rect 23716 1604 23734 1638
rect 23784 1604 23806 1638
rect 23852 1604 23878 1638
rect 23920 1604 23950 1638
rect 23988 1604 24022 1638
rect 24056 1604 24090 1638
rect 24128 1604 24158 1638
rect 24200 1604 24226 1638
rect 24272 1604 24294 1638
rect 22248 1548 22282 1562
rect 22248 1477 22282 1486
rect 22424 1448 22438 1482
rect 22492 1448 22510 1482
rect 22560 1448 22582 1482
rect 22628 1448 22654 1482
rect 22696 1448 22726 1482
rect 22764 1448 22798 1482
rect 22832 1448 22866 1482
rect 22904 1448 22934 1482
rect 22976 1448 23002 1482
rect 23048 1448 23070 1482
rect 23120 1448 23138 1482
rect 23192 1448 23206 1482
rect 23264 1448 23274 1482
rect 23336 1448 23342 1482
rect 23408 1448 23410 1482
rect 23444 1448 23446 1482
rect 23512 1448 23518 1482
rect 23580 1448 23590 1482
rect 23648 1448 23662 1482
rect 23716 1448 23734 1482
rect 23784 1448 23806 1482
rect 23852 1448 23878 1482
rect 23920 1448 23950 1482
rect 23988 1448 24022 1482
rect 24056 1448 24090 1482
rect 24128 1448 24158 1482
rect 24200 1448 24226 1482
rect 24272 1448 24294 1482
rect 22248 1406 22282 1410
rect 22248 1368 22282 1372
rect 22248 1292 22282 1301
rect 22424 1292 22438 1326
rect 22492 1292 22510 1326
rect 22560 1292 22582 1326
rect 22628 1292 22654 1326
rect 22696 1292 22726 1326
rect 22764 1292 22798 1326
rect 22832 1292 22866 1326
rect 22904 1292 22934 1326
rect 22976 1292 23002 1326
rect 23048 1292 23070 1326
rect 23120 1292 23138 1326
rect 23192 1292 23206 1326
rect 23264 1292 23274 1326
rect 23336 1292 23342 1326
rect 23408 1292 23410 1326
rect 23444 1292 23446 1326
rect 23512 1292 23518 1326
rect 23580 1292 23590 1326
rect 23648 1292 23662 1326
rect 23716 1292 23734 1326
rect 23784 1292 23806 1326
rect 23852 1292 23878 1326
rect 23920 1292 23950 1326
rect 23988 1292 24022 1326
rect 24056 1292 24090 1326
rect 24128 1292 24158 1326
rect 24200 1292 24226 1326
rect 24272 1292 24294 1326
rect 6379 1226 6383 1260
rect 6429 1226 6455 1260
rect 6497 1226 6527 1260
rect 6565 1226 6599 1260
rect 6633 1226 6667 1260
rect 6705 1226 6735 1260
rect 6777 1226 6803 1260
rect 6849 1226 6871 1260
rect 6921 1226 6939 1260
rect 6993 1226 7007 1260
rect 7065 1226 7075 1260
rect 7137 1226 7143 1260
rect 7209 1226 7211 1260
rect 7245 1226 7247 1260
rect 7313 1226 7319 1260
rect 7381 1226 7391 1260
rect 7449 1226 7463 1260
rect 7517 1226 7535 1260
rect 7585 1226 7607 1260
rect 7653 1226 7679 1260
rect 7721 1226 7751 1260
rect 7789 1226 7823 1260
rect 7857 1226 7891 1260
rect 7929 1226 7959 1260
rect 8001 1226 8027 1260
rect 8073 1226 8095 1260
rect 8145 1226 8163 1260
rect 8217 1226 8231 1260
rect 8289 1226 8299 1260
rect 8361 1226 8367 1260
rect 8433 1226 8435 1260
rect 8469 1226 8471 1260
rect 8537 1226 8543 1260
rect 8605 1226 8615 1260
rect 8673 1226 8687 1260
rect 8741 1226 8759 1260
rect 8809 1226 8831 1260
rect 8877 1226 8903 1260
rect 8945 1226 8975 1260
rect 9013 1226 9047 1260
rect 9081 1226 9115 1260
rect 9153 1226 9183 1260
rect 9225 1226 9251 1260
rect 9297 1226 9319 1260
rect 9529 1226 9533 1260
rect 9579 1226 9605 1260
rect 9647 1226 9677 1260
rect 9715 1226 9749 1260
rect 9783 1226 9817 1260
rect 9855 1226 9885 1260
rect 9927 1226 9953 1260
rect 9999 1226 10021 1260
rect 10071 1226 10089 1260
rect 10143 1226 10157 1260
rect 10215 1226 10225 1260
rect 10287 1226 10293 1260
rect 10359 1226 10361 1260
rect 10395 1226 10397 1260
rect 10463 1226 10469 1260
rect 10531 1226 10541 1260
rect 10599 1226 10613 1260
rect 10667 1226 10685 1260
rect 10735 1226 10757 1260
rect 10803 1226 10829 1260
rect 10871 1226 10901 1260
rect 10939 1226 10973 1260
rect 11007 1226 11041 1260
rect 11079 1226 11109 1260
rect 11151 1226 11177 1260
rect 11223 1226 11245 1260
rect 11295 1226 11313 1260
rect 11367 1226 11381 1260
rect 11439 1226 11449 1260
rect 11511 1226 11517 1260
rect 11583 1226 11585 1260
rect 11619 1226 11621 1260
rect 11687 1226 11693 1260
rect 11755 1226 11765 1260
rect 11823 1226 11837 1260
rect 11891 1226 11909 1260
rect 11959 1226 11981 1260
rect 12027 1226 12053 1260
rect 12095 1226 12125 1260
rect 12163 1226 12197 1260
rect 12231 1226 12265 1260
rect 12303 1226 12333 1260
rect 12375 1226 12401 1260
rect 12447 1226 12469 1260
rect 12679 1226 12683 1260
rect 12729 1226 12755 1260
rect 12797 1226 12827 1260
rect 12865 1226 12899 1260
rect 12933 1226 12967 1260
rect 13005 1226 13035 1260
rect 13077 1226 13103 1260
rect 13149 1226 13171 1260
rect 13221 1226 13239 1260
rect 13293 1226 13307 1260
rect 13365 1226 13375 1260
rect 13437 1226 13443 1260
rect 13509 1226 13511 1260
rect 13545 1226 13547 1260
rect 13613 1226 13619 1260
rect 13681 1226 13691 1260
rect 13749 1226 13763 1260
rect 13817 1226 13835 1260
rect 13885 1226 13907 1260
rect 13953 1226 13979 1260
rect 14021 1226 14051 1260
rect 14089 1226 14123 1260
rect 14157 1226 14191 1260
rect 14229 1226 14259 1260
rect 14301 1226 14327 1260
rect 14373 1226 14395 1260
rect 14445 1226 14463 1260
rect 14517 1226 14531 1260
rect 14589 1226 14599 1260
rect 14661 1226 14667 1260
rect 14733 1226 14735 1260
rect 14769 1226 14771 1260
rect 14837 1226 14843 1260
rect 14905 1226 14915 1260
rect 14973 1226 14987 1260
rect 15041 1226 15059 1260
rect 15109 1226 15131 1260
rect 15177 1226 15203 1260
rect 15245 1226 15275 1260
rect 15313 1226 15347 1260
rect 15381 1226 15415 1260
rect 15453 1226 15483 1260
rect 15525 1226 15551 1260
rect 15597 1226 15619 1260
rect 15829 1226 15833 1260
rect 15879 1226 15905 1260
rect 15947 1226 15977 1260
rect 16015 1226 16049 1260
rect 16083 1226 16117 1260
rect 16155 1226 16185 1260
rect 16227 1226 16253 1260
rect 16299 1226 16321 1260
rect 16371 1226 16389 1260
rect 16443 1226 16457 1260
rect 16515 1226 16525 1260
rect 16587 1226 16593 1260
rect 16659 1226 16661 1260
rect 16695 1226 16697 1260
rect 16763 1226 16769 1260
rect 16831 1226 16841 1260
rect 16899 1226 16913 1260
rect 16967 1226 16985 1260
rect 17035 1226 17057 1260
rect 17103 1226 17129 1260
rect 17171 1226 17201 1260
rect 17239 1226 17273 1260
rect 17307 1226 17341 1260
rect 17379 1226 17409 1260
rect 17451 1226 17477 1260
rect 17523 1226 17545 1260
rect 17595 1226 17613 1260
rect 17667 1226 17681 1260
rect 17739 1226 17749 1260
rect 17811 1226 17817 1260
rect 17883 1226 17885 1260
rect 17919 1226 17921 1260
rect 17987 1226 17993 1260
rect 18055 1226 18065 1260
rect 18123 1226 18137 1260
rect 18191 1226 18209 1260
rect 18259 1226 18281 1260
rect 18327 1226 18353 1260
rect 18395 1226 18425 1260
rect 18463 1226 18497 1260
rect 18531 1226 18565 1260
rect 18603 1226 18633 1260
rect 18675 1226 18701 1260
rect 18747 1226 18769 1260
rect 18979 1226 18983 1260
rect 19029 1226 19055 1260
rect 19097 1226 19127 1260
rect 19165 1226 19199 1260
rect 19233 1226 19267 1260
rect 19305 1226 19335 1260
rect 19377 1226 19403 1260
rect 19449 1226 19471 1260
rect 19521 1226 19539 1260
rect 19593 1226 19607 1260
rect 19665 1226 19675 1260
rect 19737 1226 19743 1260
rect 19809 1226 19811 1260
rect 19845 1226 19847 1260
rect 19913 1226 19919 1260
rect 19981 1226 19991 1260
rect 20049 1226 20063 1260
rect 20117 1226 20135 1260
rect 20185 1226 20207 1260
rect 20253 1226 20279 1260
rect 20321 1226 20351 1260
rect 20389 1226 20423 1260
rect 20457 1226 20491 1260
rect 20529 1226 20559 1260
rect 20601 1226 20627 1260
rect 20673 1226 20695 1260
rect 20745 1226 20763 1260
rect 20817 1226 20831 1260
rect 20889 1226 20899 1260
rect 20961 1226 20967 1260
rect 21033 1226 21035 1260
rect 21069 1226 21071 1260
rect 21137 1226 21143 1260
rect 21205 1226 21215 1260
rect 21273 1226 21287 1260
rect 21341 1226 21359 1260
rect 21409 1226 21431 1260
rect 21477 1226 21503 1260
rect 21545 1226 21575 1260
rect 21613 1226 21647 1260
rect 21681 1226 21715 1260
rect 21753 1226 21783 1260
rect 21825 1226 21851 1260
rect 21897 1226 21919 1260
rect 22248 1216 22282 1230
rect 6256 1193 6339 1209
rect 6256 1143 6273 1193
rect 6307 1143 6339 1193
rect 9404 1199 9489 1215
rect 9404 1183 9423 1199
rect 9422 1165 9423 1183
rect 9457 1183 9489 1199
rect 12553 1199 12639 1215
rect 12553 1183 12573 1199
rect 9457 1165 9460 1183
rect 9422 1149 9460 1165
rect 12572 1165 12573 1183
rect 12607 1183 12639 1199
rect 15703 1199 15789 1215
rect 15703 1183 15723 1199
rect 12607 1165 12610 1183
rect 12572 1149 12610 1165
rect 15722 1165 15723 1183
rect 15757 1183 15789 1199
rect 18853 1199 18939 1215
rect 18853 1183 18873 1199
rect 15757 1165 15760 1183
rect 15722 1149 15760 1165
rect 18872 1165 18873 1183
rect 18907 1183 18939 1199
rect 22003 1199 22089 1215
rect 22003 1183 22023 1199
rect 18907 1165 18910 1183
rect 18872 1149 18910 1165
rect 22022 1165 22023 1183
rect 22057 1183 22089 1199
rect 22057 1165 22060 1183
rect 22022 1149 22060 1165
rect 6256 1115 6339 1143
rect 6256 1068 6273 1115
rect 6307 1068 6339 1115
rect 9404 1128 9489 1149
rect 6379 1070 6383 1104
rect 6429 1070 6455 1104
rect 6497 1070 6527 1104
rect 6565 1070 6599 1104
rect 6633 1070 6667 1104
rect 6705 1070 6735 1104
rect 6777 1070 6803 1104
rect 6849 1070 6871 1104
rect 6921 1070 6939 1104
rect 6993 1070 7007 1104
rect 7065 1070 7075 1104
rect 7137 1070 7143 1104
rect 7209 1070 7211 1104
rect 7245 1070 7247 1104
rect 7313 1070 7319 1104
rect 7381 1070 7391 1104
rect 7449 1070 7463 1104
rect 7517 1070 7535 1104
rect 7585 1070 7607 1104
rect 7653 1070 7679 1104
rect 7721 1070 7751 1104
rect 7789 1070 7823 1104
rect 7857 1070 7891 1104
rect 7929 1070 7959 1104
rect 8001 1070 8027 1104
rect 8073 1070 8095 1104
rect 8145 1070 8163 1104
rect 8217 1070 8231 1104
rect 8289 1070 8299 1104
rect 8361 1070 8367 1104
rect 8433 1070 8435 1104
rect 8469 1070 8471 1104
rect 8537 1070 8543 1104
rect 8605 1070 8615 1104
rect 8673 1070 8687 1104
rect 8741 1070 8759 1104
rect 8809 1070 8831 1104
rect 8877 1070 8903 1104
rect 8945 1070 8975 1104
rect 9013 1070 9047 1104
rect 9081 1070 9115 1104
rect 9153 1070 9183 1104
rect 9225 1070 9251 1104
rect 9297 1070 9319 1104
rect 9404 1094 9423 1128
rect 9457 1094 9489 1128
rect 12553 1128 12639 1149
rect 6256 1037 6339 1068
rect 6256 993 6273 1037
rect 6307 993 6339 1037
rect 9404 1057 9489 1094
rect 9529 1070 9533 1104
rect 9579 1070 9605 1104
rect 9647 1070 9677 1104
rect 9715 1070 9749 1104
rect 9783 1070 9817 1104
rect 9855 1070 9885 1104
rect 9927 1070 9953 1104
rect 9999 1070 10021 1104
rect 10071 1070 10089 1104
rect 10143 1070 10157 1104
rect 10215 1070 10225 1104
rect 10287 1070 10293 1104
rect 10359 1070 10361 1104
rect 10395 1070 10397 1104
rect 10463 1070 10469 1104
rect 10531 1070 10541 1104
rect 10599 1070 10613 1104
rect 10667 1070 10685 1104
rect 10735 1070 10757 1104
rect 10803 1070 10829 1104
rect 10871 1070 10901 1104
rect 10939 1070 10973 1104
rect 11007 1070 11041 1104
rect 11079 1070 11109 1104
rect 11151 1070 11177 1104
rect 11223 1070 11245 1104
rect 11295 1070 11313 1104
rect 11367 1070 11381 1104
rect 11439 1070 11449 1104
rect 11511 1070 11517 1104
rect 11583 1070 11585 1104
rect 11619 1070 11621 1104
rect 11687 1070 11693 1104
rect 11755 1070 11765 1104
rect 11823 1070 11837 1104
rect 11891 1070 11909 1104
rect 11959 1070 11981 1104
rect 12027 1070 12053 1104
rect 12095 1070 12125 1104
rect 12163 1070 12197 1104
rect 12231 1070 12265 1104
rect 12303 1070 12333 1104
rect 12375 1070 12401 1104
rect 12447 1070 12469 1104
rect 12553 1094 12573 1128
rect 12607 1094 12639 1128
rect 15703 1128 15789 1149
rect 9404 1027 9423 1057
rect 9422 1023 9423 1027
rect 9457 1027 9489 1057
rect 12553 1057 12639 1094
rect 12679 1070 12683 1104
rect 12729 1070 12755 1104
rect 12797 1070 12827 1104
rect 12865 1070 12899 1104
rect 12933 1070 12967 1104
rect 13005 1070 13035 1104
rect 13077 1070 13103 1104
rect 13149 1070 13171 1104
rect 13221 1070 13239 1104
rect 13293 1070 13307 1104
rect 13365 1070 13375 1104
rect 13437 1070 13443 1104
rect 13509 1070 13511 1104
rect 13545 1070 13547 1104
rect 13613 1070 13619 1104
rect 13681 1070 13691 1104
rect 13749 1070 13763 1104
rect 13817 1070 13835 1104
rect 13885 1070 13907 1104
rect 13953 1070 13979 1104
rect 14021 1070 14051 1104
rect 14089 1070 14123 1104
rect 14157 1070 14191 1104
rect 14229 1070 14259 1104
rect 14301 1070 14327 1104
rect 14373 1070 14395 1104
rect 14445 1070 14463 1104
rect 14517 1070 14531 1104
rect 14589 1070 14599 1104
rect 14661 1070 14667 1104
rect 14733 1070 14735 1104
rect 14769 1070 14771 1104
rect 14837 1070 14843 1104
rect 14905 1070 14915 1104
rect 14973 1070 14987 1104
rect 15041 1070 15059 1104
rect 15109 1070 15131 1104
rect 15177 1070 15203 1104
rect 15245 1070 15275 1104
rect 15313 1070 15347 1104
rect 15381 1070 15415 1104
rect 15453 1070 15483 1104
rect 15525 1070 15551 1104
rect 15597 1070 15619 1104
rect 15703 1094 15723 1128
rect 15757 1094 15789 1128
rect 18853 1128 18939 1149
rect 12553 1027 12573 1057
rect 9457 1023 9460 1027
rect 9422 993 9460 1023
rect 12572 1023 12573 1027
rect 12607 1027 12639 1057
rect 15703 1057 15789 1094
rect 15829 1070 15833 1104
rect 15879 1070 15905 1104
rect 15947 1070 15977 1104
rect 16015 1070 16049 1104
rect 16083 1070 16117 1104
rect 16155 1070 16185 1104
rect 16227 1070 16253 1104
rect 16299 1070 16321 1104
rect 16371 1070 16389 1104
rect 16443 1070 16457 1104
rect 16515 1070 16525 1104
rect 16587 1070 16593 1104
rect 16659 1070 16661 1104
rect 16695 1070 16697 1104
rect 16763 1070 16769 1104
rect 16831 1070 16841 1104
rect 16899 1070 16913 1104
rect 16967 1070 16985 1104
rect 17035 1070 17057 1104
rect 17103 1070 17129 1104
rect 17171 1070 17201 1104
rect 17239 1070 17273 1104
rect 17307 1070 17341 1104
rect 17379 1070 17409 1104
rect 17451 1070 17477 1104
rect 17523 1070 17545 1104
rect 17595 1070 17613 1104
rect 17667 1070 17681 1104
rect 17739 1070 17749 1104
rect 17811 1070 17817 1104
rect 17883 1070 17885 1104
rect 17919 1070 17921 1104
rect 17987 1070 17993 1104
rect 18055 1070 18065 1104
rect 18123 1070 18137 1104
rect 18191 1070 18209 1104
rect 18259 1070 18281 1104
rect 18327 1070 18353 1104
rect 18395 1070 18425 1104
rect 18463 1070 18497 1104
rect 18531 1070 18565 1104
rect 18603 1070 18633 1104
rect 18675 1070 18701 1104
rect 18747 1070 18769 1104
rect 18853 1094 18873 1128
rect 18907 1094 18939 1128
rect 22003 1128 22089 1149
rect 15703 1027 15723 1057
rect 12607 1023 12610 1027
rect 12572 993 12610 1023
rect 15722 1023 15723 1027
rect 15757 1027 15789 1057
rect 18853 1057 18939 1094
rect 18979 1070 18983 1104
rect 19029 1070 19055 1104
rect 19097 1070 19127 1104
rect 19165 1070 19199 1104
rect 19233 1070 19267 1104
rect 19305 1070 19335 1104
rect 19377 1070 19403 1104
rect 19449 1070 19471 1104
rect 19521 1070 19539 1104
rect 19593 1070 19607 1104
rect 19665 1070 19675 1104
rect 19737 1070 19743 1104
rect 19809 1070 19811 1104
rect 19845 1070 19847 1104
rect 19913 1070 19919 1104
rect 19981 1070 19991 1104
rect 20049 1070 20063 1104
rect 20117 1070 20135 1104
rect 20185 1070 20207 1104
rect 20253 1070 20279 1104
rect 20321 1070 20351 1104
rect 20389 1070 20423 1104
rect 20457 1070 20491 1104
rect 20529 1070 20559 1104
rect 20601 1070 20627 1104
rect 20673 1070 20695 1104
rect 20745 1070 20763 1104
rect 20817 1070 20831 1104
rect 20889 1070 20899 1104
rect 20961 1070 20967 1104
rect 21033 1070 21035 1104
rect 21069 1070 21071 1104
rect 21137 1070 21143 1104
rect 21205 1070 21215 1104
rect 21273 1070 21287 1104
rect 21341 1070 21359 1104
rect 21409 1070 21431 1104
rect 21477 1070 21503 1104
rect 21545 1070 21575 1104
rect 21613 1070 21647 1104
rect 21681 1070 21715 1104
rect 21753 1070 21783 1104
rect 21825 1070 21851 1104
rect 21897 1070 21919 1104
rect 22003 1094 22023 1128
rect 22057 1094 22089 1128
rect 18853 1027 18873 1057
rect 15757 1023 15760 1027
rect 15722 993 15760 1023
rect 18872 1023 18873 1027
rect 18907 1027 18939 1057
rect 22003 1057 22089 1094
rect 22003 1027 22023 1057
rect 18907 1023 18910 1027
rect 18872 993 18910 1023
rect 22022 1023 22023 1027
rect 22057 1027 22089 1057
rect 22248 1140 22282 1159
rect 22424 1136 22438 1170
rect 22492 1136 22510 1170
rect 22560 1136 22582 1170
rect 22628 1136 22654 1170
rect 22696 1136 22726 1170
rect 22764 1136 22798 1170
rect 22832 1136 22866 1170
rect 22904 1136 22934 1170
rect 22976 1136 23002 1170
rect 23048 1136 23070 1170
rect 23120 1136 23138 1170
rect 23192 1136 23206 1170
rect 23264 1136 23274 1170
rect 23336 1136 23342 1170
rect 23408 1136 23410 1170
rect 23444 1136 23446 1170
rect 23512 1136 23518 1170
rect 23580 1136 23590 1170
rect 23648 1136 23662 1170
rect 23716 1136 23734 1170
rect 23784 1136 23806 1170
rect 23852 1136 23878 1170
rect 23920 1136 23950 1170
rect 23988 1136 24022 1170
rect 24056 1136 24090 1170
rect 24128 1136 24158 1170
rect 24200 1136 24226 1170
rect 24272 1136 24294 1170
rect 22248 1064 22282 1088
rect 22057 1023 22060 1027
rect 22022 993 22060 1023
rect 6256 959 6339 993
rect 6256 918 6273 959
rect 6307 918 6339 959
rect 9404 985 9489 993
rect 9404 951 9423 985
rect 9457 951 9489 985
rect 6256 881 6339 918
rect 6379 914 6383 948
rect 6429 914 6455 948
rect 6497 914 6527 948
rect 6565 914 6599 948
rect 6633 914 6667 948
rect 6705 914 6735 948
rect 6777 914 6803 948
rect 6849 914 6871 948
rect 6921 914 6939 948
rect 6993 914 7007 948
rect 7065 914 7075 948
rect 7137 914 7143 948
rect 7209 914 7211 948
rect 7245 914 7247 948
rect 7313 914 7319 948
rect 7381 914 7391 948
rect 7449 914 7463 948
rect 7517 914 7535 948
rect 7585 914 7607 948
rect 7653 914 7679 948
rect 7721 914 7751 948
rect 7789 914 7823 948
rect 7857 914 7891 948
rect 7929 914 7959 948
rect 8001 914 8027 948
rect 8073 914 8095 948
rect 8145 914 8163 948
rect 8217 914 8231 948
rect 8289 914 8299 948
rect 8361 914 8367 948
rect 8433 914 8435 948
rect 8469 914 8471 948
rect 8537 914 8543 948
rect 8605 914 8615 948
rect 8673 914 8687 948
rect 8741 914 8759 948
rect 8809 914 8831 948
rect 8877 914 8903 948
rect 8945 914 8975 948
rect 9013 914 9047 948
rect 9081 914 9115 948
rect 9153 914 9183 948
rect 9225 914 9251 948
rect 9297 914 9319 948
rect 6256 843 6273 881
rect 6307 843 6339 881
rect 9404 913 9489 951
rect 12553 985 12639 993
rect 12553 951 12573 985
rect 12607 951 12639 985
rect 9529 914 9533 948
rect 9579 914 9605 948
rect 9647 914 9677 948
rect 9715 914 9749 948
rect 9783 914 9817 948
rect 9855 914 9885 948
rect 9927 914 9953 948
rect 9999 914 10021 948
rect 10071 914 10089 948
rect 10143 914 10157 948
rect 10215 914 10225 948
rect 10287 914 10293 948
rect 10359 914 10361 948
rect 10395 914 10397 948
rect 10463 914 10469 948
rect 10531 914 10541 948
rect 10599 914 10613 948
rect 10667 914 10685 948
rect 10735 914 10757 948
rect 10803 914 10829 948
rect 10871 914 10901 948
rect 10939 914 10973 948
rect 11007 914 11041 948
rect 11079 914 11109 948
rect 11151 914 11177 948
rect 11223 914 11245 948
rect 11295 914 11313 948
rect 11367 914 11381 948
rect 11439 914 11449 948
rect 11511 914 11517 948
rect 11583 914 11585 948
rect 11619 914 11621 948
rect 11687 914 11693 948
rect 11755 914 11765 948
rect 11823 914 11837 948
rect 11891 914 11909 948
rect 11959 914 11981 948
rect 12027 914 12053 948
rect 12095 914 12125 948
rect 12163 914 12197 948
rect 12231 914 12265 948
rect 12303 914 12333 948
rect 12375 914 12401 948
rect 12447 914 12469 948
rect 9404 879 9423 913
rect 9457 879 9489 913
rect 9404 871 9489 879
rect 12553 913 12639 951
rect 15703 985 15789 993
rect 15703 951 15723 985
rect 15757 951 15789 985
rect 12679 914 12683 948
rect 12729 914 12755 948
rect 12797 914 12827 948
rect 12865 914 12899 948
rect 12933 914 12967 948
rect 13005 914 13035 948
rect 13077 914 13103 948
rect 13149 914 13171 948
rect 13221 914 13239 948
rect 13293 914 13307 948
rect 13365 914 13375 948
rect 13437 914 13443 948
rect 13509 914 13511 948
rect 13545 914 13547 948
rect 13613 914 13619 948
rect 13681 914 13691 948
rect 13749 914 13763 948
rect 13817 914 13835 948
rect 13885 914 13907 948
rect 13953 914 13979 948
rect 14021 914 14051 948
rect 14089 914 14123 948
rect 14157 914 14191 948
rect 14229 914 14259 948
rect 14301 914 14327 948
rect 14373 914 14395 948
rect 14445 914 14463 948
rect 14517 914 14531 948
rect 14589 914 14599 948
rect 14661 914 14667 948
rect 14733 914 14735 948
rect 14769 914 14771 948
rect 14837 914 14843 948
rect 14905 914 14915 948
rect 14973 914 14987 948
rect 15041 914 15059 948
rect 15109 914 15131 948
rect 15177 914 15203 948
rect 15245 914 15275 948
rect 15313 914 15347 948
rect 15381 914 15415 948
rect 15453 914 15483 948
rect 15525 914 15551 948
rect 15597 914 15619 948
rect 12553 879 12573 913
rect 12607 879 12639 913
rect 12553 871 12639 879
rect 15703 913 15789 951
rect 18853 985 18939 993
rect 18853 951 18873 985
rect 18907 951 18939 985
rect 15829 914 15833 948
rect 15879 914 15905 948
rect 15947 914 15977 948
rect 16015 914 16049 948
rect 16083 914 16117 948
rect 16155 914 16185 948
rect 16227 914 16253 948
rect 16299 914 16321 948
rect 16371 914 16389 948
rect 16443 914 16457 948
rect 16515 914 16525 948
rect 16587 914 16593 948
rect 16659 914 16661 948
rect 16695 914 16697 948
rect 16763 914 16769 948
rect 16831 914 16841 948
rect 16899 914 16913 948
rect 16967 914 16985 948
rect 17035 914 17057 948
rect 17103 914 17129 948
rect 17171 914 17201 948
rect 17239 914 17273 948
rect 17307 914 17341 948
rect 17379 914 17409 948
rect 17451 914 17477 948
rect 17523 914 17545 948
rect 17595 914 17613 948
rect 17667 914 17681 948
rect 17739 914 17749 948
rect 17811 914 17817 948
rect 17883 914 17885 948
rect 17919 914 17921 948
rect 17987 914 17993 948
rect 18055 914 18065 948
rect 18123 914 18137 948
rect 18191 914 18209 948
rect 18259 914 18281 948
rect 18327 914 18353 948
rect 18395 914 18425 948
rect 18463 914 18497 948
rect 18531 914 18565 948
rect 18603 914 18633 948
rect 18675 914 18701 948
rect 18747 914 18769 948
rect 15703 879 15723 913
rect 15757 879 15789 913
rect 15703 871 15789 879
rect 18853 913 18939 951
rect 22003 985 22089 993
rect 22003 951 22023 985
rect 22057 951 22089 985
rect 18979 914 18983 948
rect 19029 914 19055 948
rect 19097 914 19127 948
rect 19165 914 19199 948
rect 19233 914 19267 948
rect 19305 914 19335 948
rect 19377 914 19403 948
rect 19449 914 19471 948
rect 19521 914 19539 948
rect 19593 914 19607 948
rect 19665 914 19675 948
rect 19737 914 19743 948
rect 19809 914 19811 948
rect 19845 914 19847 948
rect 19913 914 19919 948
rect 19981 914 19991 948
rect 20049 914 20063 948
rect 20117 914 20135 948
rect 20185 914 20207 948
rect 20253 914 20279 948
rect 20321 914 20351 948
rect 20389 914 20423 948
rect 20457 914 20491 948
rect 20529 914 20559 948
rect 20601 914 20627 948
rect 20673 914 20695 948
rect 20745 914 20763 948
rect 20817 914 20831 948
rect 20889 914 20899 948
rect 20961 914 20967 948
rect 21033 914 21035 948
rect 21069 914 21071 948
rect 21137 914 21143 948
rect 21205 914 21215 948
rect 21273 914 21287 948
rect 21341 914 21359 948
rect 21409 914 21431 948
rect 21477 914 21503 948
rect 21545 914 21575 948
rect 21613 914 21647 948
rect 21681 914 21715 948
rect 21753 914 21783 948
rect 21825 914 21851 948
rect 21897 914 21919 948
rect 18853 879 18873 913
rect 18907 879 18939 913
rect 18853 871 18939 879
rect 22003 913 22089 951
rect 22003 879 22023 913
rect 22057 879 22089 913
rect 22003 871 22089 879
rect 22248 988 22282 1017
rect 22424 980 22438 1014
rect 22492 980 22510 1014
rect 22560 980 22582 1014
rect 22628 980 22654 1014
rect 22696 980 22726 1014
rect 22764 980 22798 1014
rect 22832 980 22866 1014
rect 22904 980 22934 1014
rect 22976 980 23002 1014
rect 23048 980 23070 1014
rect 23120 980 23138 1014
rect 23192 980 23206 1014
rect 23264 980 23274 1014
rect 23336 980 23342 1014
rect 23408 980 23410 1014
rect 23444 980 23446 1014
rect 23512 980 23518 1014
rect 23580 980 23590 1014
rect 23648 980 23662 1014
rect 23716 980 23734 1014
rect 23784 980 23806 1014
rect 23852 980 23878 1014
rect 23920 980 23950 1014
rect 23988 980 24022 1014
rect 24056 980 24090 1014
rect 24128 980 24158 1014
rect 24200 980 24226 1014
rect 24272 980 24294 1014
rect 22248 912 22282 945
rect 79 784 83 818
rect 129 784 155 818
rect 197 784 227 818
rect 265 784 299 818
rect 333 784 367 818
rect 405 784 435 818
rect 477 784 503 818
rect 549 784 571 818
rect 621 784 639 818
rect 693 784 707 818
rect 765 784 775 818
rect 837 784 843 818
rect 909 784 911 818
rect 945 784 947 818
rect 1013 784 1019 818
rect 1081 784 1091 818
rect 1149 784 1163 818
rect 1217 784 1235 818
rect 1285 784 1307 818
rect 1353 784 1379 818
rect 1421 784 1451 818
rect 1489 784 1523 818
rect 1557 784 1591 818
rect 1629 784 1659 818
rect 1701 784 1727 818
rect 1773 784 1795 818
rect 1845 784 1863 818
rect 1917 784 1931 818
rect 1989 784 1999 818
rect 2061 784 2067 818
rect 2133 784 2135 818
rect 2169 784 2171 818
rect 2237 784 2243 818
rect 2305 784 2315 818
rect 2373 784 2387 818
rect 2441 784 2459 818
rect 2509 784 2531 818
rect 2577 784 2603 818
rect 2645 784 2675 818
rect 2713 784 2747 818
rect 2781 784 2815 818
rect 2853 784 2883 818
rect 2925 784 2951 818
rect 2997 784 3019 818
rect 3103 794 3189 810
rect 3103 773 3123 794
rect 3102 760 3123 773
rect 3157 760 3189 794
rect 3229 784 3233 818
rect 3279 784 3305 818
rect 3347 784 3377 818
rect 3415 784 3449 818
rect 3483 784 3517 818
rect 3555 784 3585 818
rect 3627 784 3653 818
rect 3699 784 3721 818
rect 3771 784 3789 818
rect 3843 784 3857 818
rect 3915 784 3925 818
rect 3987 784 3993 818
rect 4059 784 4061 818
rect 4095 784 4097 818
rect 4163 784 4169 818
rect 4231 784 4241 818
rect 4299 784 4313 818
rect 4367 784 4385 818
rect 4435 784 4457 818
rect 4503 784 4529 818
rect 4571 784 4601 818
rect 4639 784 4673 818
rect 4707 784 4741 818
rect 4779 784 4809 818
rect 4851 784 4877 818
rect 4923 784 4945 818
rect 4995 784 5013 818
rect 5067 784 5081 818
rect 5139 784 5149 818
rect 5211 784 5217 818
rect 5283 784 5285 818
rect 5319 784 5321 818
rect 5387 784 5393 818
rect 5455 784 5465 818
rect 5523 784 5537 818
rect 5591 784 5609 818
rect 5659 784 5681 818
rect 5727 784 5753 818
rect 5795 784 5825 818
rect 5863 784 5897 818
rect 5931 784 5965 818
rect 6003 784 6033 818
rect 6075 784 6101 818
rect 6147 784 6169 818
rect 6256 802 6339 843
rect 9422 841 9460 871
rect 9422 837 9423 841
rect 3102 741 3189 760
rect 6256 767 6273 802
rect 6307 767 6339 802
rect 9404 807 9423 837
rect 9457 837 9460 841
rect 12572 841 12610 871
rect 12572 837 12573 841
rect 9457 807 9489 837
rect 3122 723 3160 741
rect 3122 707 3123 723
rect 3102 689 3123 707
rect 3157 707 3160 723
rect 6256 725 6339 767
rect 6379 758 6383 792
rect 6429 758 6455 792
rect 6497 758 6527 792
rect 6565 758 6599 792
rect 6633 758 6667 792
rect 6705 758 6735 792
rect 6777 758 6803 792
rect 6849 758 6871 792
rect 6921 758 6939 792
rect 6993 758 7007 792
rect 7065 758 7075 792
rect 7137 758 7143 792
rect 7209 758 7211 792
rect 7245 758 7247 792
rect 7313 758 7319 792
rect 7381 758 7391 792
rect 7449 758 7463 792
rect 7517 758 7535 792
rect 7585 758 7607 792
rect 7653 758 7679 792
rect 7721 758 7751 792
rect 7789 758 7823 792
rect 7857 758 7891 792
rect 7929 758 7959 792
rect 8001 758 8027 792
rect 8073 758 8095 792
rect 8145 758 8163 792
rect 8217 758 8231 792
rect 8289 758 8299 792
rect 8361 758 8367 792
rect 8433 758 8435 792
rect 8469 758 8471 792
rect 8537 758 8543 792
rect 8605 758 8615 792
rect 8673 758 8687 792
rect 8741 758 8759 792
rect 8809 758 8831 792
rect 8877 758 8903 792
rect 8945 758 8975 792
rect 9013 758 9047 792
rect 9081 758 9115 792
rect 9153 758 9183 792
rect 9225 758 9251 792
rect 9297 758 9319 792
rect 9404 769 9489 807
rect 12553 807 12573 837
rect 12607 837 12610 841
rect 15722 841 15760 871
rect 15722 837 15723 841
rect 12607 807 12639 837
rect 3157 689 3189 707
rect 3102 673 3189 689
rect 6256 689 6273 725
rect 6307 689 6339 725
rect 9404 735 9423 769
rect 9457 735 9489 769
rect 9529 758 9533 792
rect 9579 758 9605 792
rect 9647 758 9677 792
rect 9715 758 9749 792
rect 9783 758 9817 792
rect 9855 758 9885 792
rect 9927 758 9953 792
rect 9999 758 10021 792
rect 10071 758 10089 792
rect 10143 758 10157 792
rect 10215 758 10225 792
rect 10287 758 10293 792
rect 10359 758 10361 792
rect 10395 758 10397 792
rect 10463 758 10469 792
rect 10531 758 10541 792
rect 10599 758 10613 792
rect 10667 758 10685 792
rect 10735 758 10757 792
rect 10803 758 10829 792
rect 10871 758 10901 792
rect 10939 758 10973 792
rect 11007 758 11041 792
rect 11079 758 11109 792
rect 11151 758 11177 792
rect 11223 758 11245 792
rect 11295 758 11313 792
rect 11367 758 11381 792
rect 11439 758 11449 792
rect 11511 758 11517 792
rect 11583 758 11585 792
rect 11619 758 11621 792
rect 11687 758 11693 792
rect 11755 758 11765 792
rect 11823 758 11837 792
rect 11891 758 11909 792
rect 11959 758 11981 792
rect 12027 758 12053 792
rect 12095 758 12125 792
rect 12163 758 12197 792
rect 12231 758 12265 792
rect 12303 758 12333 792
rect 12375 758 12401 792
rect 12447 758 12469 792
rect 12553 769 12639 807
rect 15703 807 15723 837
rect 15757 837 15760 841
rect 18872 841 18910 871
rect 18872 837 18873 841
rect 15757 807 15789 837
rect 9404 715 9489 735
rect 12553 735 12573 769
rect 12607 735 12639 769
rect 12679 758 12683 792
rect 12729 758 12755 792
rect 12797 758 12827 792
rect 12865 758 12899 792
rect 12933 758 12967 792
rect 13005 758 13035 792
rect 13077 758 13103 792
rect 13149 758 13171 792
rect 13221 758 13239 792
rect 13293 758 13307 792
rect 13365 758 13375 792
rect 13437 758 13443 792
rect 13509 758 13511 792
rect 13545 758 13547 792
rect 13613 758 13619 792
rect 13681 758 13691 792
rect 13749 758 13763 792
rect 13817 758 13835 792
rect 13885 758 13907 792
rect 13953 758 13979 792
rect 14021 758 14051 792
rect 14089 758 14123 792
rect 14157 758 14191 792
rect 14229 758 14259 792
rect 14301 758 14327 792
rect 14373 758 14395 792
rect 14445 758 14463 792
rect 14517 758 14531 792
rect 14589 758 14599 792
rect 14661 758 14667 792
rect 14733 758 14735 792
rect 14769 758 14771 792
rect 14837 758 14843 792
rect 14905 758 14915 792
rect 14973 758 14987 792
rect 15041 758 15059 792
rect 15109 758 15131 792
rect 15177 758 15203 792
rect 15245 758 15275 792
rect 15313 758 15347 792
rect 15381 758 15415 792
rect 15453 758 15483 792
rect 15525 758 15551 792
rect 15597 758 15619 792
rect 15703 769 15789 807
rect 18853 807 18873 837
rect 18907 837 18910 841
rect 22022 841 22060 871
rect 22022 837 22023 841
rect 18907 807 18939 837
rect 12553 715 12639 735
rect 15703 735 15723 769
rect 15757 735 15789 769
rect 15829 758 15833 792
rect 15879 758 15905 792
rect 15947 758 15977 792
rect 16015 758 16049 792
rect 16083 758 16117 792
rect 16155 758 16185 792
rect 16227 758 16253 792
rect 16299 758 16321 792
rect 16371 758 16389 792
rect 16443 758 16457 792
rect 16515 758 16525 792
rect 16587 758 16593 792
rect 16659 758 16661 792
rect 16695 758 16697 792
rect 16763 758 16769 792
rect 16831 758 16841 792
rect 16899 758 16913 792
rect 16967 758 16985 792
rect 17035 758 17057 792
rect 17103 758 17129 792
rect 17171 758 17201 792
rect 17239 758 17273 792
rect 17307 758 17341 792
rect 17379 758 17409 792
rect 17451 758 17477 792
rect 17523 758 17545 792
rect 17595 758 17613 792
rect 17667 758 17681 792
rect 17739 758 17749 792
rect 17811 758 17817 792
rect 17883 758 17885 792
rect 17919 758 17921 792
rect 17987 758 17993 792
rect 18055 758 18065 792
rect 18123 758 18137 792
rect 18191 758 18209 792
rect 18259 758 18281 792
rect 18327 758 18353 792
rect 18395 758 18425 792
rect 18463 758 18497 792
rect 18531 758 18565 792
rect 18603 758 18633 792
rect 18675 758 18701 792
rect 18747 758 18769 792
rect 18853 769 18939 807
rect 22003 807 22023 837
rect 22057 837 22060 841
rect 22057 807 22089 837
rect 15703 715 15789 735
rect 18853 735 18873 769
rect 18907 735 18939 769
rect 18979 758 18983 792
rect 19029 758 19055 792
rect 19097 758 19127 792
rect 19165 758 19199 792
rect 19233 758 19267 792
rect 19305 758 19335 792
rect 19377 758 19403 792
rect 19449 758 19471 792
rect 19521 758 19539 792
rect 19593 758 19607 792
rect 19665 758 19675 792
rect 19737 758 19743 792
rect 19809 758 19811 792
rect 19845 758 19847 792
rect 19913 758 19919 792
rect 19981 758 19991 792
rect 20049 758 20063 792
rect 20117 758 20135 792
rect 20185 758 20207 792
rect 20253 758 20279 792
rect 20321 758 20351 792
rect 20389 758 20423 792
rect 20457 758 20491 792
rect 20529 758 20559 792
rect 20601 758 20627 792
rect 20673 758 20695 792
rect 20745 758 20763 792
rect 20817 758 20831 792
rect 20889 758 20899 792
rect 20961 758 20967 792
rect 21033 758 21035 792
rect 21069 758 21071 792
rect 21137 758 21143 792
rect 21205 758 21215 792
rect 21273 758 21287 792
rect 21341 758 21359 792
rect 21409 758 21431 792
rect 21477 758 21503 792
rect 21545 758 21575 792
rect 21613 758 21647 792
rect 21681 758 21715 792
rect 21753 758 21783 792
rect 21825 758 21851 792
rect 21897 758 21919 792
rect 22003 769 22089 807
rect 18853 715 18939 735
rect 22003 735 22023 769
rect 22057 735 22089 769
rect 22003 715 22089 735
rect 22248 836 22282 873
rect 22424 824 22438 858
rect 22492 824 22510 858
rect 22560 824 22582 858
rect 22628 824 22654 858
rect 22696 824 22726 858
rect 22764 824 22798 858
rect 22832 824 22866 858
rect 22904 824 22934 858
rect 22976 824 23002 858
rect 23048 824 23070 858
rect 23120 824 23138 858
rect 23192 824 23206 858
rect 23264 824 23274 858
rect 23336 824 23342 858
rect 23408 824 23410 858
rect 23444 824 23446 858
rect 23512 824 23518 858
rect 23580 824 23590 858
rect 23648 824 23662 858
rect 23716 824 23734 858
rect 23784 824 23806 858
rect 23852 824 23878 858
rect 23920 824 23950 858
rect 23988 824 24022 858
rect 24056 824 24090 858
rect 24128 824 24158 858
rect 24200 824 24226 858
rect 24272 824 24294 858
rect 22248 763 22282 801
rect 79 628 83 662
rect 129 628 155 662
rect 197 628 227 662
rect 265 628 299 662
rect 333 628 367 662
rect 405 628 435 662
rect 477 628 503 662
rect 549 628 571 662
rect 621 628 639 662
rect 693 628 707 662
rect 765 628 775 662
rect 837 628 843 662
rect 909 628 911 662
rect 945 628 947 662
rect 1013 628 1019 662
rect 1081 628 1091 662
rect 1149 628 1163 662
rect 1217 628 1235 662
rect 1285 628 1307 662
rect 1353 628 1379 662
rect 1421 628 1451 662
rect 1489 628 1523 662
rect 1557 628 1591 662
rect 1629 628 1659 662
rect 1701 628 1727 662
rect 1773 628 1795 662
rect 1845 628 1863 662
rect 1917 628 1931 662
rect 1989 628 1999 662
rect 2061 628 2067 662
rect 2133 628 2135 662
rect 2169 628 2171 662
rect 2237 628 2243 662
rect 2305 628 2315 662
rect 2373 628 2387 662
rect 2441 628 2459 662
rect 2509 628 2531 662
rect 2577 628 2603 662
rect 2645 628 2675 662
rect 2713 628 2747 662
rect 2781 628 2815 662
rect 2853 628 2883 662
rect 2925 628 2951 662
rect 2997 628 3019 662
rect 3229 628 3233 662
rect 3279 628 3305 662
rect 3347 628 3377 662
rect 3415 628 3449 662
rect 3483 628 3517 662
rect 3555 628 3585 662
rect 3627 628 3653 662
rect 3699 628 3721 662
rect 3771 628 3789 662
rect 3843 628 3857 662
rect 3915 628 3925 662
rect 3987 628 3993 662
rect 4059 628 4061 662
rect 4095 628 4097 662
rect 4163 628 4169 662
rect 4231 628 4241 662
rect 4299 628 4313 662
rect 4367 628 4385 662
rect 4435 628 4457 662
rect 4503 628 4529 662
rect 4571 628 4601 662
rect 4639 628 4673 662
rect 4707 628 4741 662
rect 4779 628 4809 662
rect 4851 628 4877 662
rect 4923 628 4945 662
rect 4995 628 5013 662
rect 5067 628 5081 662
rect 5139 628 5149 662
rect 5211 628 5217 662
rect 5283 628 5285 662
rect 5319 628 5321 662
rect 5387 628 5393 662
rect 5455 628 5465 662
rect 5523 628 5537 662
rect 5591 628 5609 662
rect 5659 628 5681 662
rect 5727 628 5753 662
rect 5795 628 5825 662
rect 5863 628 5897 662
rect 5931 628 5965 662
rect 6003 628 6033 662
rect 6075 628 6101 662
rect 6147 628 6169 662
rect 6256 647 6339 689
rect 9422 697 9460 715
rect 9422 681 9423 697
rect 9404 663 9423 681
rect 9457 681 9460 697
rect 12572 697 12610 715
rect 12572 681 12573 697
rect 9457 663 9489 681
rect 9404 647 9489 663
rect 12553 663 12573 681
rect 12607 681 12610 697
rect 15722 697 15760 715
rect 15722 681 15723 697
rect 12607 663 12639 681
rect 12553 647 12639 663
rect 15703 663 15723 681
rect 15757 681 15760 697
rect 18872 697 18910 715
rect 18872 681 18873 697
rect 15757 663 15789 681
rect 15703 647 15789 663
rect 18853 663 18873 681
rect 18907 681 18910 697
rect 22022 697 22060 715
rect 22022 681 22023 697
rect 18907 663 18939 681
rect 18853 647 18939 663
rect 22003 663 22023 681
rect 22057 681 22060 697
rect 22248 713 22282 726
rect 22057 663 22089 681
rect 22424 668 22438 702
rect 22492 668 22510 702
rect 22560 668 22582 702
rect 22628 668 22654 702
rect 22696 668 22726 702
rect 22764 668 22798 702
rect 22832 668 22866 702
rect 22904 668 22934 702
rect 22976 668 23002 702
rect 23048 668 23070 702
rect 23120 668 23138 702
rect 23192 668 23206 702
rect 23264 668 23274 702
rect 23336 668 23342 702
rect 23408 668 23410 702
rect 23444 668 23446 702
rect 23512 668 23518 702
rect 23580 668 23590 702
rect 23648 668 23662 702
rect 23716 668 23734 702
rect 23784 668 23806 702
rect 23852 668 23878 702
rect 23920 668 23950 702
rect 23988 668 24022 702
rect 24056 668 24090 702
rect 24128 668 24158 702
rect 24200 668 24226 702
rect 24272 668 24294 702
rect 22003 647 22089 663
rect 6379 602 6383 636
rect 6429 602 6455 636
rect 6497 602 6527 636
rect 6565 602 6599 636
rect 6633 602 6667 636
rect 6705 602 6735 636
rect 6777 602 6803 636
rect 6849 602 6871 636
rect 6921 602 6939 636
rect 6993 602 7007 636
rect 7065 602 7075 636
rect 7137 602 7143 636
rect 7209 602 7211 636
rect 7245 602 7247 636
rect 7313 602 7319 636
rect 7381 602 7391 636
rect 7449 602 7463 636
rect 7517 602 7535 636
rect 7585 602 7607 636
rect 7653 602 7679 636
rect 7721 602 7751 636
rect 7789 602 7823 636
rect 7857 602 7891 636
rect 7929 602 7959 636
rect 8001 602 8027 636
rect 8073 602 8095 636
rect 8145 602 8163 636
rect 8217 602 8231 636
rect 8289 602 8299 636
rect 8361 602 8367 636
rect 8433 602 8435 636
rect 8469 602 8471 636
rect 8537 602 8543 636
rect 8605 602 8615 636
rect 8673 602 8687 636
rect 8741 602 8759 636
rect 8809 602 8831 636
rect 8877 602 8903 636
rect 8945 602 8975 636
rect 9013 602 9047 636
rect 9081 602 9115 636
rect 9153 602 9183 636
rect 9225 602 9251 636
rect 9297 602 9319 636
rect 9529 602 9533 636
rect 9579 602 9605 636
rect 9647 602 9677 636
rect 9715 602 9749 636
rect 9783 602 9817 636
rect 9855 602 9885 636
rect 9927 602 9953 636
rect 9999 602 10021 636
rect 10071 602 10089 636
rect 10143 602 10157 636
rect 10215 602 10225 636
rect 10287 602 10293 636
rect 10359 602 10361 636
rect 10395 602 10397 636
rect 10463 602 10469 636
rect 10531 602 10541 636
rect 10599 602 10613 636
rect 10667 602 10685 636
rect 10735 602 10757 636
rect 10803 602 10829 636
rect 10871 602 10901 636
rect 10939 602 10973 636
rect 11007 602 11041 636
rect 11079 602 11109 636
rect 11151 602 11177 636
rect 11223 602 11245 636
rect 11295 602 11313 636
rect 11367 602 11381 636
rect 11439 602 11449 636
rect 11511 602 11517 636
rect 11583 602 11585 636
rect 11619 602 11621 636
rect 11687 602 11693 636
rect 11755 602 11765 636
rect 11823 602 11837 636
rect 11891 602 11909 636
rect 11959 602 11981 636
rect 12027 602 12053 636
rect 12095 602 12125 636
rect 12163 602 12197 636
rect 12231 602 12265 636
rect 12303 602 12333 636
rect 12375 602 12401 636
rect 12447 602 12469 636
rect 12679 602 12683 636
rect 12729 602 12755 636
rect 12797 602 12827 636
rect 12865 602 12899 636
rect 12933 602 12967 636
rect 13005 602 13035 636
rect 13077 602 13103 636
rect 13149 602 13171 636
rect 13221 602 13239 636
rect 13293 602 13307 636
rect 13365 602 13375 636
rect 13437 602 13443 636
rect 13509 602 13511 636
rect 13545 602 13547 636
rect 13613 602 13619 636
rect 13681 602 13691 636
rect 13749 602 13763 636
rect 13817 602 13835 636
rect 13885 602 13907 636
rect 13953 602 13979 636
rect 14021 602 14051 636
rect 14089 602 14123 636
rect 14157 602 14191 636
rect 14229 602 14259 636
rect 14301 602 14327 636
rect 14373 602 14395 636
rect 14445 602 14463 636
rect 14517 602 14531 636
rect 14589 602 14599 636
rect 14661 602 14667 636
rect 14733 602 14735 636
rect 14769 602 14771 636
rect 14837 602 14843 636
rect 14905 602 14915 636
rect 14973 602 14987 636
rect 15041 602 15059 636
rect 15109 602 15131 636
rect 15177 602 15203 636
rect 15245 602 15275 636
rect 15313 602 15347 636
rect 15381 602 15415 636
rect 15453 602 15483 636
rect 15525 602 15551 636
rect 15597 602 15619 636
rect 15829 602 15833 636
rect 15879 602 15905 636
rect 15947 602 15977 636
rect 16015 602 16049 636
rect 16083 602 16117 636
rect 16155 602 16185 636
rect 16227 602 16253 636
rect 16299 602 16321 636
rect 16371 602 16389 636
rect 16443 602 16457 636
rect 16515 602 16525 636
rect 16587 602 16593 636
rect 16659 602 16661 636
rect 16695 602 16697 636
rect 16763 602 16769 636
rect 16831 602 16841 636
rect 16899 602 16913 636
rect 16967 602 16985 636
rect 17035 602 17057 636
rect 17103 602 17129 636
rect 17171 602 17201 636
rect 17239 602 17273 636
rect 17307 602 17341 636
rect 17379 602 17409 636
rect 17451 602 17477 636
rect 17523 602 17545 636
rect 17595 602 17613 636
rect 17667 602 17681 636
rect 17739 602 17749 636
rect 17811 602 17817 636
rect 17883 602 17885 636
rect 17919 602 17921 636
rect 17987 602 17993 636
rect 18055 602 18065 636
rect 18123 602 18137 636
rect 18191 602 18209 636
rect 18259 602 18281 636
rect 18327 602 18353 636
rect 18395 602 18425 636
rect 18463 602 18497 636
rect 18531 602 18565 636
rect 18603 602 18633 636
rect 18675 602 18701 636
rect 18747 602 18769 636
rect 18979 602 18983 636
rect 19029 602 19055 636
rect 19097 602 19127 636
rect 19165 602 19199 636
rect 19233 602 19267 636
rect 19305 602 19335 636
rect 19377 602 19403 636
rect 19449 602 19471 636
rect 19521 602 19539 636
rect 19593 602 19607 636
rect 19665 602 19675 636
rect 19737 602 19743 636
rect 19809 602 19811 636
rect 19845 602 19847 636
rect 19913 602 19919 636
rect 19981 602 19991 636
rect 20049 602 20063 636
rect 20117 602 20135 636
rect 20185 602 20207 636
rect 20253 602 20279 636
rect 20321 602 20351 636
rect 20389 602 20423 636
rect 20457 602 20491 636
rect 20529 602 20559 636
rect 20601 602 20627 636
rect 20673 602 20695 636
rect 20745 602 20763 636
rect 20817 602 20831 636
rect 20889 602 20899 636
rect 20961 602 20967 636
rect 21033 602 21035 636
rect 21069 602 21071 636
rect 21137 602 21143 636
rect 21205 602 21215 636
rect 21273 602 21287 636
rect 21341 602 21359 636
rect 21409 602 21431 636
rect 21477 602 21503 636
rect 21545 602 21575 636
rect 21613 602 21647 636
rect 21681 602 21715 636
rect 21753 602 21783 636
rect 21825 602 21851 636
rect 21897 602 21919 636
<< viali >>
rect 22366 2072 22390 2106
rect 22390 2072 22400 2106
rect 22438 2072 22458 2106
rect 22458 2072 22472 2106
rect 22510 2072 22526 2106
rect 22526 2072 22544 2106
rect 22582 2072 22594 2106
rect 22594 2072 22616 2106
rect 22654 2072 22662 2106
rect 22662 2072 22688 2106
rect 22726 2072 22730 2106
rect 22730 2072 22760 2106
rect 22798 2072 22832 2106
rect 22870 2072 22900 2106
rect 22900 2072 22904 2106
rect 22942 2072 22968 2106
rect 22968 2072 22976 2106
rect 23014 2072 23036 2106
rect 23036 2072 23048 2106
rect 23086 2072 23104 2106
rect 23104 2072 23120 2106
rect 23158 2072 23172 2106
rect 23172 2072 23192 2106
rect 23230 2072 23240 2106
rect 23240 2072 23264 2106
rect 23302 2072 23308 2106
rect 23308 2072 23336 2106
rect 23374 2072 23376 2106
rect 23376 2072 23408 2106
rect 23446 2072 23478 2106
rect 23478 2072 23480 2106
rect 23518 2072 23546 2106
rect 23546 2072 23552 2106
rect 23590 2072 23614 2106
rect 23614 2072 23624 2106
rect 23662 2072 23682 2106
rect 23682 2072 23696 2106
rect 23734 2072 23750 2106
rect 23750 2072 23768 2106
rect 23806 2072 23818 2106
rect 23818 2072 23840 2106
rect 23878 2072 23886 2106
rect 23886 2072 23912 2106
rect 23950 2072 23954 2106
rect 23954 2072 23984 2106
rect 24022 2072 24056 2106
rect 24094 2072 24124 2106
rect 24124 2072 24128 2106
rect 24166 2072 24192 2106
rect 24192 2072 24200 2106
rect 24238 2072 24260 2106
rect 24260 2072 24272 2106
rect 24310 2072 24328 2106
rect 24328 2072 24344 2106
rect 22248 2045 22282 2049
rect 22248 2015 22282 2045
rect 22248 1940 22282 1974
rect 22366 1916 22390 1950
rect 22390 1916 22400 1950
rect 22438 1916 22458 1950
rect 22458 1916 22472 1950
rect 22510 1916 22526 1950
rect 22526 1916 22544 1950
rect 22582 1916 22594 1950
rect 22594 1916 22616 1950
rect 22654 1916 22662 1950
rect 22662 1916 22688 1950
rect 22726 1916 22730 1950
rect 22730 1916 22760 1950
rect 22798 1916 22832 1950
rect 22870 1916 22900 1950
rect 22900 1916 22904 1950
rect 22942 1916 22968 1950
rect 22968 1916 22976 1950
rect 23014 1916 23036 1950
rect 23036 1916 23048 1950
rect 23086 1916 23104 1950
rect 23104 1916 23120 1950
rect 23158 1916 23172 1950
rect 23172 1916 23192 1950
rect 23230 1916 23240 1950
rect 23240 1916 23264 1950
rect 23302 1916 23308 1950
rect 23308 1916 23336 1950
rect 23374 1916 23376 1950
rect 23376 1916 23408 1950
rect 23446 1916 23478 1950
rect 23478 1916 23480 1950
rect 23518 1916 23546 1950
rect 23546 1916 23552 1950
rect 23590 1916 23614 1950
rect 23614 1916 23624 1950
rect 23662 1916 23682 1950
rect 23682 1916 23696 1950
rect 23734 1916 23750 1950
rect 23750 1916 23768 1950
rect 23806 1916 23818 1950
rect 23818 1916 23840 1950
rect 23878 1916 23886 1950
rect 23886 1916 23912 1950
rect 23950 1916 23954 1950
rect 23954 1916 23984 1950
rect 24022 1916 24056 1950
rect 24094 1916 24124 1950
rect 24124 1916 24128 1950
rect 24166 1916 24192 1950
rect 24192 1916 24200 1950
rect 24238 1916 24260 1950
rect 24260 1916 24272 1950
rect 24310 1916 24328 1950
rect 24328 1916 24344 1950
rect 22248 1869 22282 1899
rect 22248 1865 22282 1869
rect 22248 1798 22282 1824
rect 22248 1790 22282 1798
rect 22366 1760 22390 1794
rect 22390 1760 22400 1794
rect 22438 1760 22458 1794
rect 22458 1760 22472 1794
rect 22510 1760 22526 1794
rect 22526 1760 22544 1794
rect 22582 1760 22594 1794
rect 22594 1760 22616 1794
rect 22654 1760 22662 1794
rect 22662 1760 22688 1794
rect 22726 1760 22730 1794
rect 22730 1760 22760 1794
rect 22798 1760 22832 1794
rect 22870 1760 22900 1794
rect 22900 1760 22904 1794
rect 22942 1760 22968 1794
rect 22968 1760 22976 1794
rect 23014 1760 23036 1794
rect 23036 1760 23048 1794
rect 23086 1760 23104 1794
rect 23104 1760 23120 1794
rect 23158 1760 23172 1794
rect 23172 1760 23192 1794
rect 23230 1760 23240 1794
rect 23240 1760 23264 1794
rect 23302 1760 23308 1794
rect 23308 1760 23336 1794
rect 23374 1760 23376 1794
rect 23376 1760 23408 1794
rect 23446 1760 23478 1794
rect 23478 1760 23480 1794
rect 23518 1760 23546 1794
rect 23546 1760 23552 1794
rect 23590 1760 23614 1794
rect 23614 1760 23624 1794
rect 23662 1760 23682 1794
rect 23682 1760 23696 1794
rect 23734 1760 23750 1794
rect 23750 1760 23768 1794
rect 23806 1760 23818 1794
rect 23818 1760 23840 1794
rect 23878 1760 23886 1794
rect 23886 1760 23912 1794
rect 23950 1760 23954 1794
rect 23954 1760 23984 1794
rect 24022 1760 24056 1794
rect 24094 1760 24124 1794
rect 24124 1760 24128 1794
rect 24166 1760 24192 1794
rect 24192 1760 24200 1794
rect 24238 1760 24260 1794
rect 24260 1760 24272 1794
rect 24310 1760 24328 1794
rect 24328 1760 24344 1794
rect 22248 1727 22282 1748
rect 22248 1714 22282 1727
rect 22248 1656 22282 1672
rect 22248 1638 22282 1656
rect 22366 1604 22390 1638
rect 22390 1604 22400 1638
rect 22438 1604 22458 1638
rect 22458 1604 22472 1638
rect 22510 1604 22526 1638
rect 22526 1604 22544 1638
rect 22582 1604 22594 1638
rect 22594 1604 22616 1638
rect 22654 1604 22662 1638
rect 22662 1604 22688 1638
rect 22726 1604 22730 1638
rect 22730 1604 22760 1638
rect 22798 1604 22832 1638
rect 22870 1604 22900 1638
rect 22900 1604 22904 1638
rect 22942 1604 22968 1638
rect 22968 1604 22976 1638
rect 23014 1604 23036 1638
rect 23036 1604 23048 1638
rect 23086 1604 23104 1638
rect 23104 1604 23120 1638
rect 23158 1604 23172 1638
rect 23172 1604 23192 1638
rect 23230 1604 23240 1638
rect 23240 1604 23264 1638
rect 23302 1604 23308 1638
rect 23308 1604 23336 1638
rect 23374 1604 23376 1638
rect 23376 1604 23408 1638
rect 23446 1604 23478 1638
rect 23478 1604 23480 1638
rect 23518 1604 23546 1638
rect 23546 1604 23552 1638
rect 23590 1604 23614 1638
rect 23614 1604 23624 1638
rect 23662 1604 23682 1638
rect 23682 1604 23696 1638
rect 23734 1604 23750 1638
rect 23750 1604 23768 1638
rect 23806 1604 23818 1638
rect 23818 1604 23840 1638
rect 23878 1604 23886 1638
rect 23886 1604 23912 1638
rect 23950 1604 23954 1638
rect 23954 1604 23984 1638
rect 24022 1604 24056 1638
rect 24094 1604 24124 1638
rect 24124 1604 24128 1638
rect 24166 1604 24192 1638
rect 24192 1604 24200 1638
rect 24238 1604 24260 1638
rect 24260 1604 24272 1638
rect 24310 1604 24328 1638
rect 24328 1604 24344 1638
rect 22248 1585 22282 1596
rect 22248 1562 22282 1585
rect 22248 1514 22282 1520
rect 22248 1486 22282 1514
rect 22366 1448 22390 1482
rect 22390 1448 22400 1482
rect 22438 1448 22458 1482
rect 22458 1448 22472 1482
rect 22510 1448 22526 1482
rect 22526 1448 22544 1482
rect 22582 1448 22594 1482
rect 22594 1448 22616 1482
rect 22654 1448 22662 1482
rect 22662 1448 22688 1482
rect 22726 1448 22730 1482
rect 22730 1448 22760 1482
rect 22798 1448 22832 1482
rect 22870 1448 22900 1482
rect 22900 1448 22904 1482
rect 22942 1448 22968 1482
rect 22968 1448 22976 1482
rect 23014 1448 23036 1482
rect 23036 1448 23048 1482
rect 23086 1448 23104 1482
rect 23104 1448 23120 1482
rect 23158 1448 23172 1482
rect 23172 1448 23192 1482
rect 23230 1448 23240 1482
rect 23240 1448 23264 1482
rect 23302 1448 23308 1482
rect 23308 1448 23336 1482
rect 23374 1448 23376 1482
rect 23376 1448 23408 1482
rect 23446 1448 23478 1482
rect 23478 1448 23480 1482
rect 23518 1448 23546 1482
rect 23546 1448 23552 1482
rect 23590 1448 23614 1482
rect 23614 1448 23624 1482
rect 23662 1448 23682 1482
rect 23682 1448 23696 1482
rect 23734 1448 23750 1482
rect 23750 1448 23768 1482
rect 23806 1448 23818 1482
rect 23818 1448 23840 1482
rect 23878 1448 23886 1482
rect 23886 1448 23912 1482
rect 23950 1448 23954 1482
rect 23954 1448 23984 1482
rect 24022 1448 24056 1482
rect 24094 1448 24124 1482
rect 24124 1448 24128 1482
rect 24166 1448 24192 1482
rect 24192 1448 24200 1482
rect 24238 1448 24260 1482
rect 24260 1448 24272 1482
rect 24310 1448 24328 1482
rect 24328 1448 24344 1482
rect 22248 1443 22282 1444
rect 22248 1410 22282 1443
rect 22248 1335 22282 1368
rect 22248 1334 22282 1335
rect 22366 1292 22390 1326
rect 22390 1292 22400 1326
rect 22438 1292 22458 1326
rect 22458 1292 22472 1326
rect 22510 1292 22526 1326
rect 22526 1292 22544 1326
rect 22582 1292 22594 1326
rect 22594 1292 22616 1326
rect 22654 1292 22662 1326
rect 22662 1292 22688 1326
rect 22726 1292 22730 1326
rect 22730 1292 22760 1326
rect 22798 1292 22832 1326
rect 22870 1292 22900 1326
rect 22900 1292 22904 1326
rect 22942 1292 22968 1326
rect 22968 1292 22976 1326
rect 23014 1292 23036 1326
rect 23036 1292 23048 1326
rect 23086 1292 23104 1326
rect 23104 1292 23120 1326
rect 23158 1292 23172 1326
rect 23172 1292 23192 1326
rect 23230 1292 23240 1326
rect 23240 1292 23264 1326
rect 23302 1292 23308 1326
rect 23308 1292 23336 1326
rect 23374 1292 23376 1326
rect 23376 1292 23408 1326
rect 23446 1292 23478 1326
rect 23478 1292 23480 1326
rect 23518 1292 23546 1326
rect 23546 1292 23552 1326
rect 23590 1292 23614 1326
rect 23614 1292 23624 1326
rect 23662 1292 23682 1326
rect 23682 1292 23696 1326
rect 23734 1292 23750 1326
rect 23750 1292 23768 1326
rect 23806 1292 23818 1326
rect 23818 1292 23840 1326
rect 23878 1292 23886 1326
rect 23886 1292 23912 1326
rect 23950 1292 23954 1326
rect 23954 1292 23984 1326
rect 24022 1292 24056 1326
rect 24094 1292 24124 1326
rect 24124 1292 24128 1326
rect 24166 1292 24192 1326
rect 24192 1292 24200 1326
rect 24238 1292 24260 1326
rect 24260 1292 24272 1326
rect 24310 1292 24328 1326
rect 24328 1292 24344 1326
rect 22248 1264 22282 1292
rect 6383 1226 6395 1260
rect 6395 1226 6417 1260
rect 6455 1226 6463 1260
rect 6463 1226 6489 1260
rect 6527 1226 6531 1260
rect 6531 1226 6561 1260
rect 6599 1226 6633 1260
rect 6671 1226 6701 1260
rect 6701 1226 6705 1260
rect 6743 1226 6769 1260
rect 6769 1226 6777 1260
rect 6815 1226 6837 1260
rect 6837 1226 6849 1260
rect 6887 1226 6905 1260
rect 6905 1226 6921 1260
rect 6959 1226 6973 1260
rect 6973 1226 6993 1260
rect 7031 1226 7041 1260
rect 7041 1226 7065 1260
rect 7103 1226 7109 1260
rect 7109 1226 7137 1260
rect 7175 1226 7177 1260
rect 7177 1226 7209 1260
rect 7247 1226 7279 1260
rect 7279 1226 7281 1260
rect 7319 1226 7347 1260
rect 7347 1226 7353 1260
rect 7391 1226 7415 1260
rect 7415 1226 7425 1260
rect 7463 1226 7483 1260
rect 7483 1226 7497 1260
rect 7535 1226 7551 1260
rect 7551 1226 7569 1260
rect 7607 1226 7619 1260
rect 7619 1226 7641 1260
rect 7679 1226 7687 1260
rect 7687 1226 7713 1260
rect 7751 1226 7755 1260
rect 7755 1226 7785 1260
rect 7823 1226 7857 1260
rect 7895 1226 7925 1260
rect 7925 1226 7929 1260
rect 7967 1226 7993 1260
rect 7993 1226 8001 1260
rect 8039 1226 8061 1260
rect 8061 1226 8073 1260
rect 8111 1226 8129 1260
rect 8129 1226 8145 1260
rect 8183 1226 8197 1260
rect 8197 1226 8217 1260
rect 8255 1226 8265 1260
rect 8265 1226 8289 1260
rect 8327 1226 8333 1260
rect 8333 1226 8361 1260
rect 8399 1226 8401 1260
rect 8401 1226 8433 1260
rect 8471 1226 8503 1260
rect 8503 1226 8505 1260
rect 8543 1226 8571 1260
rect 8571 1226 8577 1260
rect 8615 1226 8639 1260
rect 8639 1226 8649 1260
rect 8687 1226 8707 1260
rect 8707 1226 8721 1260
rect 8759 1226 8775 1260
rect 8775 1226 8793 1260
rect 8831 1226 8843 1260
rect 8843 1226 8865 1260
rect 8903 1226 8911 1260
rect 8911 1226 8937 1260
rect 8975 1226 8979 1260
rect 8979 1226 9009 1260
rect 9047 1226 9081 1260
rect 9119 1226 9149 1260
rect 9149 1226 9153 1260
rect 9191 1226 9217 1260
rect 9217 1226 9225 1260
rect 9263 1226 9285 1260
rect 9285 1226 9297 1260
rect 9335 1226 9353 1260
rect 9353 1226 9369 1260
rect 9533 1226 9545 1260
rect 9545 1226 9567 1260
rect 9605 1226 9613 1260
rect 9613 1226 9639 1260
rect 9677 1226 9681 1260
rect 9681 1226 9711 1260
rect 9749 1226 9783 1260
rect 9821 1226 9851 1260
rect 9851 1226 9855 1260
rect 9893 1226 9919 1260
rect 9919 1226 9927 1260
rect 9965 1226 9987 1260
rect 9987 1226 9999 1260
rect 10037 1226 10055 1260
rect 10055 1226 10071 1260
rect 10109 1226 10123 1260
rect 10123 1226 10143 1260
rect 10181 1226 10191 1260
rect 10191 1226 10215 1260
rect 10253 1226 10259 1260
rect 10259 1226 10287 1260
rect 10325 1226 10327 1260
rect 10327 1226 10359 1260
rect 10397 1226 10429 1260
rect 10429 1226 10431 1260
rect 10469 1226 10497 1260
rect 10497 1226 10503 1260
rect 10541 1226 10565 1260
rect 10565 1226 10575 1260
rect 10613 1226 10633 1260
rect 10633 1226 10647 1260
rect 10685 1226 10701 1260
rect 10701 1226 10719 1260
rect 10757 1226 10769 1260
rect 10769 1226 10791 1260
rect 10829 1226 10837 1260
rect 10837 1226 10863 1260
rect 10901 1226 10905 1260
rect 10905 1226 10935 1260
rect 10973 1226 11007 1260
rect 11045 1226 11075 1260
rect 11075 1226 11079 1260
rect 11117 1226 11143 1260
rect 11143 1226 11151 1260
rect 11189 1226 11211 1260
rect 11211 1226 11223 1260
rect 11261 1226 11279 1260
rect 11279 1226 11295 1260
rect 11333 1226 11347 1260
rect 11347 1226 11367 1260
rect 11405 1226 11415 1260
rect 11415 1226 11439 1260
rect 11477 1226 11483 1260
rect 11483 1226 11511 1260
rect 11549 1226 11551 1260
rect 11551 1226 11583 1260
rect 11621 1226 11653 1260
rect 11653 1226 11655 1260
rect 11693 1226 11721 1260
rect 11721 1226 11727 1260
rect 11765 1226 11789 1260
rect 11789 1226 11799 1260
rect 11837 1226 11857 1260
rect 11857 1226 11871 1260
rect 11909 1226 11925 1260
rect 11925 1226 11943 1260
rect 11981 1226 11993 1260
rect 11993 1226 12015 1260
rect 12053 1226 12061 1260
rect 12061 1226 12087 1260
rect 12125 1226 12129 1260
rect 12129 1226 12159 1260
rect 12197 1226 12231 1260
rect 12269 1226 12299 1260
rect 12299 1226 12303 1260
rect 12341 1226 12367 1260
rect 12367 1226 12375 1260
rect 12413 1226 12435 1260
rect 12435 1226 12447 1260
rect 12485 1226 12503 1260
rect 12503 1226 12519 1260
rect 12683 1226 12695 1260
rect 12695 1226 12717 1260
rect 12755 1226 12763 1260
rect 12763 1226 12789 1260
rect 12827 1226 12831 1260
rect 12831 1226 12861 1260
rect 12899 1226 12933 1260
rect 12971 1226 13001 1260
rect 13001 1226 13005 1260
rect 13043 1226 13069 1260
rect 13069 1226 13077 1260
rect 13115 1226 13137 1260
rect 13137 1226 13149 1260
rect 13187 1226 13205 1260
rect 13205 1226 13221 1260
rect 13259 1226 13273 1260
rect 13273 1226 13293 1260
rect 13331 1226 13341 1260
rect 13341 1226 13365 1260
rect 13403 1226 13409 1260
rect 13409 1226 13437 1260
rect 13475 1226 13477 1260
rect 13477 1226 13509 1260
rect 13547 1226 13579 1260
rect 13579 1226 13581 1260
rect 13619 1226 13647 1260
rect 13647 1226 13653 1260
rect 13691 1226 13715 1260
rect 13715 1226 13725 1260
rect 13763 1226 13783 1260
rect 13783 1226 13797 1260
rect 13835 1226 13851 1260
rect 13851 1226 13869 1260
rect 13907 1226 13919 1260
rect 13919 1226 13941 1260
rect 13979 1226 13987 1260
rect 13987 1226 14013 1260
rect 14051 1226 14055 1260
rect 14055 1226 14085 1260
rect 14123 1226 14157 1260
rect 14195 1226 14225 1260
rect 14225 1226 14229 1260
rect 14267 1226 14293 1260
rect 14293 1226 14301 1260
rect 14339 1226 14361 1260
rect 14361 1226 14373 1260
rect 14411 1226 14429 1260
rect 14429 1226 14445 1260
rect 14483 1226 14497 1260
rect 14497 1226 14517 1260
rect 14555 1226 14565 1260
rect 14565 1226 14589 1260
rect 14627 1226 14633 1260
rect 14633 1226 14661 1260
rect 14699 1226 14701 1260
rect 14701 1226 14733 1260
rect 14771 1226 14803 1260
rect 14803 1226 14805 1260
rect 14843 1226 14871 1260
rect 14871 1226 14877 1260
rect 14915 1226 14939 1260
rect 14939 1226 14949 1260
rect 14987 1226 15007 1260
rect 15007 1226 15021 1260
rect 15059 1226 15075 1260
rect 15075 1226 15093 1260
rect 15131 1226 15143 1260
rect 15143 1226 15165 1260
rect 15203 1226 15211 1260
rect 15211 1226 15237 1260
rect 15275 1226 15279 1260
rect 15279 1226 15309 1260
rect 15347 1226 15381 1260
rect 15419 1226 15449 1260
rect 15449 1226 15453 1260
rect 15491 1226 15517 1260
rect 15517 1226 15525 1260
rect 15563 1226 15585 1260
rect 15585 1226 15597 1260
rect 15635 1226 15653 1260
rect 15653 1226 15669 1260
rect 15833 1226 15845 1260
rect 15845 1226 15867 1260
rect 15905 1226 15913 1260
rect 15913 1226 15939 1260
rect 15977 1226 15981 1260
rect 15981 1226 16011 1260
rect 16049 1226 16083 1260
rect 16121 1226 16151 1260
rect 16151 1226 16155 1260
rect 16193 1226 16219 1260
rect 16219 1226 16227 1260
rect 16265 1226 16287 1260
rect 16287 1226 16299 1260
rect 16337 1226 16355 1260
rect 16355 1226 16371 1260
rect 16409 1226 16423 1260
rect 16423 1226 16443 1260
rect 16481 1226 16491 1260
rect 16491 1226 16515 1260
rect 16553 1226 16559 1260
rect 16559 1226 16587 1260
rect 16625 1226 16627 1260
rect 16627 1226 16659 1260
rect 16697 1226 16729 1260
rect 16729 1226 16731 1260
rect 16769 1226 16797 1260
rect 16797 1226 16803 1260
rect 16841 1226 16865 1260
rect 16865 1226 16875 1260
rect 16913 1226 16933 1260
rect 16933 1226 16947 1260
rect 16985 1226 17001 1260
rect 17001 1226 17019 1260
rect 17057 1226 17069 1260
rect 17069 1226 17091 1260
rect 17129 1226 17137 1260
rect 17137 1226 17163 1260
rect 17201 1226 17205 1260
rect 17205 1226 17235 1260
rect 17273 1226 17307 1260
rect 17345 1226 17375 1260
rect 17375 1226 17379 1260
rect 17417 1226 17443 1260
rect 17443 1226 17451 1260
rect 17489 1226 17511 1260
rect 17511 1226 17523 1260
rect 17561 1226 17579 1260
rect 17579 1226 17595 1260
rect 17633 1226 17647 1260
rect 17647 1226 17667 1260
rect 17705 1226 17715 1260
rect 17715 1226 17739 1260
rect 17777 1226 17783 1260
rect 17783 1226 17811 1260
rect 17849 1226 17851 1260
rect 17851 1226 17883 1260
rect 17921 1226 17953 1260
rect 17953 1226 17955 1260
rect 17993 1226 18021 1260
rect 18021 1226 18027 1260
rect 18065 1226 18089 1260
rect 18089 1226 18099 1260
rect 18137 1226 18157 1260
rect 18157 1226 18171 1260
rect 18209 1226 18225 1260
rect 18225 1226 18243 1260
rect 18281 1226 18293 1260
rect 18293 1226 18315 1260
rect 18353 1226 18361 1260
rect 18361 1226 18387 1260
rect 18425 1226 18429 1260
rect 18429 1226 18459 1260
rect 18497 1226 18531 1260
rect 18569 1226 18599 1260
rect 18599 1226 18603 1260
rect 18641 1226 18667 1260
rect 18667 1226 18675 1260
rect 18713 1226 18735 1260
rect 18735 1226 18747 1260
rect 18785 1226 18803 1260
rect 18803 1226 18819 1260
rect 18983 1226 18995 1260
rect 18995 1226 19017 1260
rect 19055 1226 19063 1260
rect 19063 1226 19089 1260
rect 19127 1226 19131 1260
rect 19131 1226 19161 1260
rect 19199 1226 19233 1260
rect 19271 1226 19301 1260
rect 19301 1226 19305 1260
rect 19343 1226 19369 1260
rect 19369 1226 19377 1260
rect 19415 1226 19437 1260
rect 19437 1226 19449 1260
rect 19487 1226 19505 1260
rect 19505 1226 19521 1260
rect 19559 1226 19573 1260
rect 19573 1226 19593 1260
rect 19631 1226 19641 1260
rect 19641 1226 19665 1260
rect 19703 1226 19709 1260
rect 19709 1226 19737 1260
rect 19775 1226 19777 1260
rect 19777 1226 19809 1260
rect 19847 1226 19879 1260
rect 19879 1226 19881 1260
rect 19919 1226 19947 1260
rect 19947 1226 19953 1260
rect 19991 1226 20015 1260
rect 20015 1226 20025 1260
rect 20063 1226 20083 1260
rect 20083 1226 20097 1260
rect 20135 1226 20151 1260
rect 20151 1226 20169 1260
rect 20207 1226 20219 1260
rect 20219 1226 20241 1260
rect 20279 1226 20287 1260
rect 20287 1226 20313 1260
rect 20351 1226 20355 1260
rect 20355 1226 20385 1260
rect 20423 1226 20457 1260
rect 20495 1226 20525 1260
rect 20525 1226 20529 1260
rect 20567 1226 20593 1260
rect 20593 1226 20601 1260
rect 20639 1226 20661 1260
rect 20661 1226 20673 1260
rect 20711 1226 20729 1260
rect 20729 1226 20745 1260
rect 20783 1226 20797 1260
rect 20797 1226 20817 1260
rect 20855 1226 20865 1260
rect 20865 1226 20889 1260
rect 20927 1226 20933 1260
rect 20933 1226 20961 1260
rect 20999 1226 21001 1260
rect 21001 1226 21033 1260
rect 21071 1226 21103 1260
rect 21103 1226 21105 1260
rect 21143 1226 21171 1260
rect 21171 1226 21177 1260
rect 21215 1226 21239 1260
rect 21239 1226 21249 1260
rect 21287 1226 21307 1260
rect 21307 1226 21321 1260
rect 21359 1226 21375 1260
rect 21375 1226 21393 1260
rect 21431 1226 21443 1260
rect 21443 1226 21465 1260
rect 21503 1226 21511 1260
rect 21511 1226 21537 1260
rect 21575 1226 21579 1260
rect 21579 1226 21609 1260
rect 21647 1226 21681 1260
rect 21719 1226 21749 1260
rect 21749 1226 21753 1260
rect 21791 1226 21817 1260
rect 21817 1226 21825 1260
rect 21863 1226 21885 1260
rect 21885 1226 21897 1260
rect 21935 1226 21953 1260
rect 21953 1226 21969 1260
rect 22248 1258 22282 1264
rect 6273 1159 6307 1177
rect 6273 1143 6307 1159
rect 9388 1149 9422 1183
rect 9460 1149 9494 1183
rect 12538 1149 12572 1183
rect 12610 1149 12644 1183
rect 15688 1149 15722 1183
rect 15760 1149 15794 1183
rect 18838 1149 18872 1183
rect 18910 1149 18944 1183
rect 21988 1149 22022 1183
rect 22248 1193 22282 1216
rect 22060 1149 22094 1183
rect 22248 1182 22282 1193
rect 6273 1081 6307 1102
rect 6273 1068 6307 1081
rect 6383 1070 6395 1104
rect 6395 1070 6417 1104
rect 6455 1070 6463 1104
rect 6463 1070 6489 1104
rect 6527 1070 6531 1104
rect 6531 1070 6561 1104
rect 6599 1070 6633 1104
rect 6671 1070 6701 1104
rect 6701 1070 6705 1104
rect 6743 1070 6769 1104
rect 6769 1070 6777 1104
rect 6815 1070 6837 1104
rect 6837 1070 6849 1104
rect 6887 1070 6905 1104
rect 6905 1070 6921 1104
rect 6959 1070 6973 1104
rect 6973 1070 6993 1104
rect 7031 1070 7041 1104
rect 7041 1070 7065 1104
rect 7103 1070 7109 1104
rect 7109 1070 7137 1104
rect 7175 1070 7177 1104
rect 7177 1070 7209 1104
rect 7247 1070 7279 1104
rect 7279 1070 7281 1104
rect 7319 1070 7347 1104
rect 7347 1070 7353 1104
rect 7391 1070 7415 1104
rect 7415 1070 7425 1104
rect 7463 1070 7483 1104
rect 7483 1070 7497 1104
rect 7535 1070 7551 1104
rect 7551 1070 7569 1104
rect 7607 1070 7619 1104
rect 7619 1070 7641 1104
rect 7679 1070 7687 1104
rect 7687 1070 7713 1104
rect 7751 1070 7755 1104
rect 7755 1070 7785 1104
rect 7823 1070 7857 1104
rect 7895 1070 7925 1104
rect 7925 1070 7929 1104
rect 7967 1070 7993 1104
rect 7993 1070 8001 1104
rect 8039 1070 8061 1104
rect 8061 1070 8073 1104
rect 8111 1070 8129 1104
rect 8129 1070 8145 1104
rect 8183 1070 8197 1104
rect 8197 1070 8217 1104
rect 8255 1070 8265 1104
rect 8265 1070 8289 1104
rect 8327 1070 8333 1104
rect 8333 1070 8361 1104
rect 8399 1070 8401 1104
rect 8401 1070 8433 1104
rect 8471 1070 8503 1104
rect 8503 1070 8505 1104
rect 8543 1070 8571 1104
rect 8571 1070 8577 1104
rect 8615 1070 8639 1104
rect 8639 1070 8649 1104
rect 8687 1070 8707 1104
rect 8707 1070 8721 1104
rect 8759 1070 8775 1104
rect 8775 1070 8793 1104
rect 8831 1070 8843 1104
rect 8843 1070 8865 1104
rect 8903 1070 8911 1104
rect 8911 1070 8937 1104
rect 8975 1070 8979 1104
rect 8979 1070 9009 1104
rect 9047 1070 9081 1104
rect 9119 1070 9149 1104
rect 9149 1070 9153 1104
rect 9191 1070 9217 1104
rect 9217 1070 9225 1104
rect 9263 1070 9285 1104
rect 9285 1070 9297 1104
rect 9335 1070 9353 1104
rect 9353 1070 9369 1104
rect 6273 1003 6307 1027
rect 6273 993 6307 1003
rect 9533 1070 9545 1104
rect 9545 1070 9567 1104
rect 9605 1070 9613 1104
rect 9613 1070 9639 1104
rect 9677 1070 9681 1104
rect 9681 1070 9711 1104
rect 9749 1070 9783 1104
rect 9821 1070 9851 1104
rect 9851 1070 9855 1104
rect 9893 1070 9919 1104
rect 9919 1070 9927 1104
rect 9965 1070 9987 1104
rect 9987 1070 9999 1104
rect 10037 1070 10055 1104
rect 10055 1070 10071 1104
rect 10109 1070 10123 1104
rect 10123 1070 10143 1104
rect 10181 1070 10191 1104
rect 10191 1070 10215 1104
rect 10253 1070 10259 1104
rect 10259 1070 10287 1104
rect 10325 1070 10327 1104
rect 10327 1070 10359 1104
rect 10397 1070 10429 1104
rect 10429 1070 10431 1104
rect 10469 1070 10497 1104
rect 10497 1070 10503 1104
rect 10541 1070 10565 1104
rect 10565 1070 10575 1104
rect 10613 1070 10633 1104
rect 10633 1070 10647 1104
rect 10685 1070 10701 1104
rect 10701 1070 10719 1104
rect 10757 1070 10769 1104
rect 10769 1070 10791 1104
rect 10829 1070 10837 1104
rect 10837 1070 10863 1104
rect 10901 1070 10905 1104
rect 10905 1070 10935 1104
rect 10973 1070 11007 1104
rect 11045 1070 11075 1104
rect 11075 1070 11079 1104
rect 11117 1070 11143 1104
rect 11143 1070 11151 1104
rect 11189 1070 11211 1104
rect 11211 1070 11223 1104
rect 11261 1070 11279 1104
rect 11279 1070 11295 1104
rect 11333 1070 11347 1104
rect 11347 1070 11367 1104
rect 11405 1070 11415 1104
rect 11415 1070 11439 1104
rect 11477 1070 11483 1104
rect 11483 1070 11511 1104
rect 11549 1070 11551 1104
rect 11551 1070 11583 1104
rect 11621 1070 11653 1104
rect 11653 1070 11655 1104
rect 11693 1070 11721 1104
rect 11721 1070 11727 1104
rect 11765 1070 11789 1104
rect 11789 1070 11799 1104
rect 11837 1070 11857 1104
rect 11857 1070 11871 1104
rect 11909 1070 11925 1104
rect 11925 1070 11943 1104
rect 11981 1070 11993 1104
rect 11993 1070 12015 1104
rect 12053 1070 12061 1104
rect 12061 1070 12087 1104
rect 12125 1070 12129 1104
rect 12129 1070 12159 1104
rect 12197 1070 12231 1104
rect 12269 1070 12299 1104
rect 12299 1070 12303 1104
rect 12341 1070 12367 1104
rect 12367 1070 12375 1104
rect 12413 1070 12435 1104
rect 12435 1070 12447 1104
rect 12485 1070 12503 1104
rect 12503 1070 12519 1104
rect 9388 993 9422 1027
rect 12683 1070 12695 1104
rect 12695 1070 12717 1104
rect 12755 1070 12763 1104
rect 12763 1070 12789 1104
rect 12827 1070 12831 1104
rect 12831 1070 12861 1104
rect 12899 1070 12933 1104
rect 12971 1070 13001 1104
rect 13001 1070 13005 1104
rect 13043 1070 13069 1104
rect 13069 1070 13077 1104
rect 13115 1070 13137 1104
rect 13137 1070 13149 1104
rect 13187 1070 13205 1104
rect 13205 1070 13221 1104
rect 13259 1070 13273 1104
rect 13273 1070 13293 1104
rect 13331 1070 13341 1104
rect 13341 1070 13365 1104
rect 13403 1070 13409 1104
rect 13409 1070 13437 1104
rect 13475 1070 13477 1104
rect 13477 1070 13509 1104
rect 13547 1070 13579 1104
rect 13579 1070 13581 1104
rect 13619 1070 13647 1104
rect 13647 1070 13653 1104
rect 13691 1070 13715 1104
rect 13715 1070 13725 1104
rect 13763 1070 13783 1104
rect 13783 1070 13797 1104
rect 13835 1070 13851 1104
rect 13851 1070 13869 1104
rect 13907 1070 13919 1104
rect 13919 1070 13941 1104
rect 13979 1070 13987 1104
rect 13987 1070 14013 1104
rect 14051 1070 14055 1104
rect 14055 1070 14085 1104
rect 14123 1070 14157 1104
rect 14195 1070 14225 1104
rect 14225 1070 14229 1104
rect 14267 1070 14293 1104
rect 14293 1070 14301 1104
rect 14339 1070 14361 1104
rect 14361 1070 14373 1104
rect 14411 1070 14429 1104
rect 14429 1070 14445 1104
rect 14483 1070 14497 1104
rect 14497 1070 14517 1104
rect 14555 1070 14565 1104
rect 14565 1070 14589 1104
rect 14627 1070 14633 1104
rect 14633 1070 14661 1104
rect 14699 1070 14701 1104
rect 14701 1070 14733 1104
rect 14771 1070 14803 1104
rect 14803 1070 14805 1104
rect 14843 1070 14871 1104
rect 14871 1070 14877 1104
rect 14915 1070 14939 1104
rect 14939 1070 14949 1104
rect 14987 1070 15007 1104
rect 15007 1070 15021 1104
rect 15059 1070 15075 1104
rect 15075 1070 15093 1104
rect 15131 1070 15143 1104
rect 15143 1070 15165 1104
rect 15203 1070 15211 1104
rect 15211 1070 15237 1104
rect 15275 1070 15279 1104
rect 15279 1070 15309 1104
rect 15347 1070 15381 1104
rect 15419 1070 15449 1104
rect 15449 1070 15453 1104
rect 15491 1070 15517 1104
rect 15517 1070 15525 1104
rect 15563 1070 15585 1104
rect 15585 1070 15597 1104
rect 15635 1070 15653 1104
rect 15653 1070 15669 1104
rect 9460 993 9494 1027
rect 12538 993 12572 1027
rect 15833 1070 15845 1104
rect 15845 1070 15867 1104
rect 15905 1070 15913 1104
rect 15913 1070 15939 1104
rect 15977 1070 15981 1104
rect 15981 1070 16011 1104
rect 16049 1070 16083 1104
rect 16121 1070 16151 1104
rect 16151 1070 16155 1104
rect 16193 1070 16219 1104
rect 16219 1070 16227 1104
rect 16265 1070 16287 1104
rect 16287 1070 16299 1104
rect 16337 1070 16355 1104
rect 16355 1070 16371 1104
rect 16409 1070 16423 1104
rect 16423 1070 16443 1104
rect 16481 1070 16491 1104
rect 16491 1070 16515 1104
rect 16553 1070 16559 1104
rect 16559 1070 16587 1104
rect 16625 1070 16627 1104
rect 16627 1070 16659 1104
rect 16697 1070 16729 1104
rect 16729 1070 16731 1104
rect 16769 1070 16797 1104
rect 16797 1070 16803 1104
rect 16841 1070 16865 1104
rect 16865 1070 16875 1104
rect 16913 1070 16933 1104
rect 16933 1070 16947 1104
rect 16985 1070 17001 1104
rect 17001 1070 17019 1104
rect 17057 1070 17069 1104
rect 17069 1070 17091 1104
rect 17129 1070 17137 1104
rect 17137 1070 17163 1104
rect 17201 1070 17205 1104
rect 17205 1070 17235 1104
rect 17273 1070 17307 1104
rect 17345 1070 17375 1104
rect 17375 1070 17379 1104
rect 17417 1070 17443 1104
rect 17443 1070 17451 1104
rect 17489 1070 17511 1104
rect 17511 1070 17523 1104
rect 17561 1070 17579 1104
rect 17579 1070 17595 1104
rect 17633 1070 17647 1104
rect 17647 1070 17667 1104
rect 17705 1070 17715 1104
rect 17715 1070 17739 1104
rect 17777 1070 17783 1104
rect 17783 1070 17811 1104
rect 17849 1070 17851 1104
rect 17851 1070 17883 1104
rect 17921 1070 17953 1104
rect 17953 1070 17955 1104
rect 17993 1070 18021 1104
rect 18021 1070 18027 1104
rect 18065 1070 18089 1104
rect 18089 1070 18099 1104
rect 18137 1070 18157 1104
rect 18157 1070 18171 1104
rect 18209 1070 18225 1104
rect 18225 1070 18243 1104
rect 18281 1070 18293 1104
rect 18293 1070 18315 1104
rect 18353 1070 18361 1104
rect 18361 1070 18387 1104
rect 18425 1070 18429 1104
rect 18429 1070 18459 1104
rect 18497 1070 18531 1104
rect 18569 1070 18599 1104
rect 18599 1070 18603 1104
rect 18641 1070 18667 1104
rect 18667 1070 18675 1104
rect 18713 1070 18735 1104
rect 18735 1070 18747 1104
rect 18785 1070 18803 1104
rect 18803 1070 18819 1104
rect 12610 993 12644 1027
rect 15688 993 15722 1027
rect 18983 1070 18995 1104
rect 18995 1070 19017 1104
rect 19055 1070 19063 1104
rect 19063 1070 19089 1104
rect 19127 1070 19131 1104
rect 19131 1070 19161 1104
rect 19199 1070 19233 1104
rect 19271 1070 19301 1104
rect 19301 1070 19305 1104
rect 19343 1070 19369 1104
rect 19369 1070 19377 1104
rect 19415 1070 19437 1104
rect 19437 1070 19449 1104
rect 19487 1070 19505 1104
rect 19505 1070 19521 1104
rect 19559 1070 19573 1104
rect 19573 1070 19593 1104
rect 19631 1070 19641 1104
rect 19641 1070 19665 1104
rect 19703 1070 19709 1104
rect 19709 1070 19737 1104
rect 19775 1070 19777 1104
rect 19777 1070 19809 1104
rect 19847 1070 19879 1104
rect 19879 1070 19881 1104
rect 19919 1070 19947 1104
rect 19947 1070 19953 1104
rect 19991 1070 20015 1104
rect 20015 1070 20025 1104
rect 20063 1070 20083 1104
rect 20083 1070 20097 1104
rect 20135 1070 20151 1104
rect 20151 1070 20169 1104
rect 20207 1070 20219 1104
rect 20219 1070 20241 1104
rect 20279 1070 20287 1104
rect 20287 1070 20313 1104
rect 20351 1070 20355 1104
rect 20355 1070 20385 1104
rect 20423 1070 20457 1104
rect 20495 1070 20525 1104
rect 20525 1070 20529 1104
rect 20567 1070 20593 1104
rect 20593 1070 20601 1104
rect 20639 1070 20661 1104
rect 20661 1070 20673 1104
rect 20711 1070 20729 1104
rect 20729 1070 20745 1104
rect 20783 1070 20797 1104
rect 20797 1070 20817 1104
rect 20855 1070 20865 1104
rect 20865 1070 20889 1104
rect 20927 1070 20933 1104
rect 20933 1070 20961 1104
rect 20999 1070 21001 1104
rect 21001 1070 21033 1104
rect 21071 1070 21103 1104
rect 21103 1070 21105 1104
rect 21143 1070 21171 1104
rect 21171 1070 21177 1104
rect 21215 1070 21239 1104
rect 21239 1070 21249 1104
rect 21287 1070 21307 1104
rect 21307 1070 21321 1104
rect 21359 1070 21375 1104
rect 21375 1070 21393 1104
rect 21431 1070 21443 1104
rect 21443 1070 21465 1104
rect 21503 1070 21511 1104
rect 21511 1070 21537 1104
rect 21575 1070 21579 1104
rect 21579 1070 21609 1104
rect 21647 1070 21681 1104
rect 21719 1070 21749 1104
rect 21749 1070 21753 1104
rect 21791 1070 21817 1104
rect 21817 1070 21825 1104
rect 21863 1070 21885 1104
rect 21885 1070 21897 1104
rect 21935 1070 21953 1104
rect 21953 1070 21969 1104
rect 15760 993 15794 1027
rect 18838 993 18872 1027
rect 18910 993 18944 1027
rect 21988 993 22022 1027
rect 22248 1122 22282 1140
rect 22366 1136 22390 1170
rect 22390 1136 22400 1170
rect 22438 1136 22458 1170
rect 22458 1136 22472 1170
rect 22510 1136 22526 1170
rect 22526 1136 22544 1170
rect 22582 1136 22594 1170
rect 22594 1136 22616 1170
rect 22654 1136 22662 1170
rect 22662 1136 22688 1170
rect 22726 1136 22730 1170
rect 22730 1136 22760 1170
rect 22798 1136 22832 1170
rect 22870 1136 22900 1170
rect 22900 1136 22904 1170
rect 22942 1136 22968 1170
rect 22968 1136 22976 1170
rect 23014 1136 23036 1170
rect 23036 1136 23048 1170
rect 23086 1136 23104 1170
rect 23104 1136 23120 1170
rect 23158 1136 23172 1170
rect 23172 1136 23192 1170
rect 23230 1136 23240 1170
rect 23240 1136 23264 1170
rect 23302 1136 23308 1170
rect 23308 1136 23336 1170
rect 23374 1136 23376 1170
rect 23376 1136 23408 1170
rect 23446 1136 23478 1170
rect 23478 1136 23480 1170
rect 23518 1136 23546 1170
rect 23546 1136 23552 1170
rect 23590 1136 23614 1170
rect 23614 1136 23624 1170
rect 23662 1136 23682 1170
rect 23682 1136 23696 1170
rect 23734 1136 23750 1170
rect 23750 1136 23768 1170
rect 23806 1136 23818 1170
rect 23818 1136 23840 1170
rect 23878 1136 23886 1170
rect 23886 1136 23912 1170
rect 23950 1136 23954 1170
rect 23954 1136 23984 1170
rect 24022 1136 24056 1170
rect 24094 1136 24124 1170
rect 24124 1136 24128 1170
rect 24166 1136 24192 1170
rect 24192 1136 24200 1170
rect 24238 1136 24260 1170
rect 24260 1136 24272 1170
rect 24310 1136 24328 1170
rect 24328 1136 24344 1170
rect 22248 1106 22282 1122
rect 22248 1051 22282 1064
rect 22248 1030 22282 1051
rect 22060 993 22094 1027
rect 6273 925 6307 952
rect 6273 918 6307 925
rect 6383 914 6395 948
rect 6395 914 6417 948
rect 6455 914 6463 948
rect 6463 914 6489 948
rect 6527 914 6531 948
rect 6531 914 6561 948
rect 6599 914 6633 948
rect 6671 914 6701 948
rect 6701 914 6705 948
rect 6743 914 6769 948
rect 6769 914 6777 948
rect 6815 914 6837 948
rect 6837 914 6849 948
rect 6887 914 6905 948
rect 6905 914 6921 948
rect 6959 914 6973 948
rect 6973 914 6993 948
rect 7031 914 7041 948
rect 7041 914 7065 948
rect 7103 914 7109 948
rect 7109 914 7137 948
rect 7175 914 7177 948
rect 7177 914 7209 948
rect 7247 914 7279 948
rect 7279 914 7281 948
rect 7319 914 7347 948
rect 7347 914 7353 948
rect 7391 914 7415 948
rect 7415 914 7425 948
rect 7463 914 7483 948
rect 7483 914 7497 948
rect 7535 914 7551 948
rect 7551 914 7569 948
rect 7607 914 7619 948
rect 7619 914 7641 948
rect 7679 914 7687 948
rect 7687 914 7713 948
rect 7751 914 7755 948
rect 7755 914 7785 948
rect 7823 914 7857 948
rect 7895 914 7925 948
rect 7925 914 7929 948
rect 7967 914 7993 948
rect 7993 914 8001 948
rect 8039 914 8061 948
rect 8061 914 8073 948
rect 8111 914 8129 948
rect 8129 914 8145 948
rect 8183 914 8197 948
rect 8197 914 8217 948
rect 8255 914 8265 948
rect 8265 914 8289 948
rect 8327 914 8333 948
rect 8333 914 8361 948
rect 8399 914 8401 948
rect 8401 914 8433 948
rect 8471 914 8503 948
rect 8503 914 8505 948
rect 8543 914 8571 948
rect 8571 914 8577 948
rect 8615 914 8639 948
rect 8639 914 8649 948
rect 8687 914 8707 948
rect 8707 914 8721 948
rect 8759 914 8775 948
rect 8775 914 8793 948
rect 8831 914 8843 948
rect 8843 914 8865 948
rect 8903 914 8911 948
rect 8911 914 8937 948
rect 8975 914 8979 948
rect 8979 914 9009 948
rect 9047 914 9081 948
rect 9119 914 9149 948
rect 9149 914 9153 948
rect 9191 914 9217 948
rect 9217 914 9225 948
rect 9263 914 9285 948
rect 9285 914 9297 948
rect 9335 914 9353 948
rect 9353 914 9369 948
rect 6273 847 6307 877
rect 6273 843 6307 847
rect 9533 914 9545 948
rect 9545 914 9567 948
rect 9605 914 9613 948
rect 9613 914 9639 948
rect 9677 914 9681 948
rect 9681 914 9711 948
rect 9749 914 9783 948
rect 9821 914 9851 948
rect 9851 914 9855 948
rect 9893 914 9919 948
rect 9919 914 9927 948
rect 9965 914 9987 948
rect 9987 914 9999 948
rect 10037 914 10055 948
rect 10055 914 10071 948
rect 10109 914 10123 948
rect 10123 914 10143 948
rect 10181 914 10191 948
rect 10191 914 10215 948
rect 10253 914 10259 948
rect 10259 914 10287 948
rect 10325 914 10327 948
rect 10327 914 10359 948
rect 10397 914 10429 948
rect 10429 914 10431 948
rect 10469 914 10497 948
rect 10497 914 10503 948
rect 10541 914 10565 948
rect 10565 914 10575 948
rect 10613 914 10633 948
rect 10633 914 10647 948
rect 10685 914 10701 948
rect 10701 914 10719 948
rect 10757 914 10769 948
rect 10769 914 10791 948
rect 10829 914 10837 948
rect 10837 914 10863 948
rect 10901 914 10905 948
rect 10905 914 10935 948
rect 10973 914 11007 948
rect 11045 914 11075 948
rect 11075 914 11079 948
rect 11117 914 11143 948
rect 11143 914 11151 948
rect 11189 914 11211 948
rect 11211 914 11223 948
rect 11261 914 11279 948
rect 11279 914 11295 948
rect 11333 914 11347 948
rect 11347 914 11367 948
rect 11405 914 11415 948
rect 11415 914 11439 948
rect 11477 914 11483 948
rect 11483 914 11511 948
rect 11549 914 11551 948
rect 11551 914 11583 948
rect 11621 914 11653 948
rect 11653 914 11655 948
rect 11693 914 11721 948
rect 11721 914 11727 948
rect 11765 914 11789 948
rect 11789 914 11799 948
rect 11837 914 11857 948
rect 11857 914 11871 948
rect 11909 914 11925 948
rect 11925 914 11943 948
rect 11981 914 11993 948
rect 11993 914 12015 948
rect 12053 914 12061 948
rect 12061 914 12087 948
rect 12125 914 12129 948
rect 12129 914 12159 948
rect 12197 914 12231 948
rect 12269 914 12299 948
rect 12299 914 12303 948
rect 12341 914 12367 948
rect 12367 914 12375 948
rect 12413 914 12435 948
rect 12435 914 12447 948
rect 12485 914 12503 948
rect 12503 914 12519 948
rect 12683 914 12695 948
rect 12695 914 12717 948
rect 12755 914 12763 948
rect 12763 914 12789 948
rect 12827 914 12831 948
rect 12831 914 12861 948
rect 12899 914 12933 948
rect 12971 914 13001 948
rect 13001 914 13005 948
rect 13043 914 13069 948
rect 13069 914 13077 948
rect 13115 914 13137 948
rect 13137 914 13149 948
rect 13187 914 13205 948
rect 13205 914 13221 948
rect 13259 914 13273 948
rect 13273 914 13293 948
rect 13331 914 13341 948
rect 13341 914 13365 948
rect 13403 914 13409 948
rect 13409 914 13437 948
rect 13475 914 13477 948
rect 13477 914 13509 948
rect 13547 914 13579 948
rect 13579 914 13581 948
rect 13619 914 13647 948
rect 13647 914 13653 948
rect 13691 914 13715 948
rect 13715 914 13725 948
rect 13763 914 13783 948
rect 13783 914 13797 948
rect 13835 914 13851 948
rect 13851 914 13869 948
rect 13907 914 13919 948
rect 13919 914 13941 948
rect 13979 914 13987 948
rect 13987 914 14013 948
rect 14051 914 14055 948
rect 14055 914 14085 948
rect 14123 914 14157 948
rect 14195 914 14225 948
rect 14225 914 14229 948
rect 14267 914 14293 948
rect 14293 914 14301 948
rect 14339 914 14361 948
rect 14361 914 14373 948
rect 14411 914 14429 948
rect 14429 914 14445 948
rect 14483 914 14497 948
rect 14497 914 14517 948
rect 14555 914 14565 948
rect 14565 914 14589 948
rect 14627 914 14633 948
rect 14633 914 14661 948
rect 14699 914 14701 948
rect 14701 914 14733 948
rect 14771 914 14803 948
rect 14803 914 14805 948
rect 14843 914 14871 948
rect 14871 914 14877 948
rect 14915 914 14939 948
rect 14939 914 14949 948
rect 14987 914 15007 948
rect 15007 914 15021 948
rect 15059 914 15075 948
rect 15075 914 15093 948
rect 15131 914 15143 948
rect 15143 914 15165 948
rect 15203 914 15211 948
rect 15211 914 15237 948
rect 15275 914 15279 948
rect 15279 914 15309 948
rect 15347 914 15381 948
rect 15419 914 15449 948
rect 15449 914 15453 948
rect 15491 914 15517 948
rect 15517 914 15525 948
rect 15563 914 15585 948
rect 15585 914 15597 948
rect 15635 914 15653 948
rect 15653 914 15669 948
rect 15833 914 15845 948
rect 15845 914 15867 948
rect 15905 914 15913 948
rect 15913 914 15939 948
rect 15977 914 15981 948
rect 15981 914 16011 948
rect 16049 914 16083 948
rect 16121 914 16151 948
rect 16151 914 16155 948
rect 16193 914 16219 948
rect 16219 914 16227 948
rect 16265 914 16287 948
rect 16287 914 16299 948
rect 16337 914 16355 948
rect 16355 914 16371 948
rect 16409 914 16423 948
rect 16423 914 16443 948
rect 16481 914 16491 948
rect 16491 914 16515 948
rect 16553 914 16559 948
rect 16559 914 16587 948
rect 16625 914 16627 948
rect 16627 914 16659 948
rect 16697 914 16729 948
rect 16729 914 16731 948
rect 16769 914 16797 948
rect 16797 914 16803 948
rect 16841 914 16865 948
rect 16865 914 16875 948
rect 16913 914 16933 948
rect 16933 914 16947 948
rect 16985 914 17001 948
rect 17001 914 17019 948
rect 17057 914 17069 948
rect 17069 914 17091 948
rect 17129 914 17137 948
rect 17137 914 17163 948
rect 17201 914 17205 948
rect 17205 914 17235 948
rect 17273 914 17307 948
rect 17345 914 17375 948
rect 17375 914 17379 948
rect 17417 914 17443 948
rect 17443 914 17451 948
rect 17489 914 17511 948
rect 17511 914 17523 948
rect 17561 914 17579 948
rect 17579 914 17595 948
rect 17633 914 17647 948
rect 17647 914 17667 948
rect 17705 914 17715 948
rect 17715 914 17739 948
rect 17777 914 17783 948
rect 17783 914 17811 948
rect 17849 914 17851 948
rect 17851 914 17883 948
rect 17921 914 17953 948
rect 17953 914 17955 948
rect 17993 914 18021 948
rect 18021 914 18027 948
rect 18065 914 18089 948
rect 18089 914 18099 948
rect 18137 914 18157 948
rect 18157 914 18171 948
rect 18209 914 18225 948
rect 18225 914 18243 948
rect 18281 914 18293 948
rect 18293 914 18315 948
rect 18353 914 18361 948
rect 18361 914 18387 948
rect 18425 914 18429 948
rect 18429 914 18459 948
rect 18497 914 18531 948
rect 18569 914 18599 948
rect 18599 914 18603 948
rect 18641 914 18667 948
rect 18667 914 18675 948
rect 18713 914 18735 948
rect 18735 914 18747 948
rect 18785 914 18803 948
rect 18803 914 18819 948
rect 18983 914 18995 948
rect 18995 914 19017 948
rect 19055 914 19063 948
rect 19063 914 19089 948
rect 19127 914 19131 948
rect 19131 914 19161 948
rect 19199 914 19233 948
rect 19271 914 19301 948
rect 19301 914 19305 948
rect 19343 914 19369 948
rect 19369 914 19377 948
rect 19415 914 19437 948
rect 19437 914 19449 948
rect 19487 914 19505 948
rect 19505 914 19521 948
rect 19559 914 19573 948
rect 19573 914 19593 948
rect 19631 914 19641 948
rect 19641 914 19665 948
rect 19703 914 19709 948
rect 19709 914 19737 948
rect 19775 914 19777 948
rect 19777 914 19809 948
rect 19847 914 19879 948
rect 19879 914 19881 948
rect 19919 914 19947 948
rect 19947 914 19953 948
rect 19991 914 20015 948
rect 20015 914 20025 948
rect 20063 914 20083 948
rect 20083 914 20097 948
rect 20135 914 20151 948
rect 20151 914 20169 948
rect 20207 914 20219 948
rect 20219 914 20241 948
rect 20279 914 20287 948
rect 20287 914 20313 948
rect 20351 914 20355 948
rect 20355 914 20385 948
rect 20423 914 20457 948
rect 20495 914 20525 948
rect 20525 914 20529 948
rect 20567 914 20593 948
rect 20593 914 20601 948
rect 20639 914 20661 948
rect 20661 914 20673 948
rect 20711 914 20729 948
rect 20729 914 20745 948
rect 20783 914 20797 948
rect 20797 914 20817 948
rect 20855 914 20865 948
rect 20865 914 20889 948
rect 20927 914 20933 948
rect 20933 914 20961 948
rect 20999 914 21001 948
rect 21001 914 21033 948
rect 21071 914 21103 948
rect 21103 914 21105 948
rect 21143 914 21171 948
rect 21171 914 21177 948
rect 21215 914 21239 948
rect 21239 914 21249 948
rect 21287 914 21307 948
rect 21307 914 21321 948
rect 21359 914 21375 948
rect 21375 914 21393 948
rect 21431 914 21443 948
rect 21443 914 21465 948
rect 21503 914 21511 948
rect 21511 914 21537 948
rect 21575 914 21579 948
rect 21579 914 21609 948
rect 21647 914 21681 948
rect 21719 914 21749 948
rect 21749 914 21753 948
rect 21791 914 21817 948
rect 21817 914 21825 948
rect 21863 914 21885 948
rect 21885 914 21897 948
rect 21935 914 21953 948
rect 21953 914 21969 948
rect 22248 979 22282 988
rect 22366 980 22390 1014
rect 22390 980 22400 1014
rect 22438 980 22458 1014
rect 22458 980 22472 1014
rect 22510 980 22526 1014
rect 22526 980 22544 1014
rect 22582 980 22594 1014
rect 22594 980 22616 1014
rect 22654 980 22662 1014
rect 22662 980 22688 1014
rect 22726 980 22730 1014
rect 22730 980 22760 1014
rect 22798 980 22832 1014
rect 22870 980 22900 1014
rect 22900 980 22904 1014
rect 22942 980 22968 1014
rect 22968 980 22976 1014
rect 23014 980 23036 1014
rect 23036 980 23048 1014
rect 23086 980 23104 1014
rect 23104 980 23120 1014
rect 23158 980 23172 1014
rect 23172 980 23192 1014
rect 23230 980 23240 1014
rect 23240 980 23264 1014
rect 23302 980 23308 1014
rect 23308 980 23336 1014
rect 23374 980 23376 1014
rect 23376 980 23408 1014
rect 23446 980 23478 1014
rect 23478 980 23480 1014
rect 23518 980 23546 1014
rect 23546 980 23552 1014
rect 23590 980 23614 1014
rect 23614 980 23624 1014
rect 23662 980 23682 1014
rect 23682 980 23696 1014
rect 23734 980 23750 1014
rect 23750 980 23768 1014
rect 23806 980 23818 1014
rect 23818 980 23840 1014
rect 23878 980 23886 1014
rect 23886 980 23912 1014
rect 23950 980 23954 1014
rect 23954 980 23984 1014
rect 24022 980 24056 1014
rect 24094 980 24124 1014
rect 24124 980 24128 1014
rect 24166 980 24192 1014
rect 24192 980 24200 1014
rect 24238 980 24260 1014
rect 24260 980 24272 1014
rect 24310 980 24328 1014
rect 24328 980 24344 1014
rect 22248 954 22282 979
rect 22248 907 22282 912
rect 22248 878 22282 907
rect 83 784 95 818
rect 95 784 117 818
rect 155 784 163 818
rect 163 784 189 818
rect 227 784 231 818
rect 231 784 261 818
rect 299 784 333 818
rect 371 784 401 818
rect 401 784 405 818
rect 443 784 469 818
rect 469 784 477 818
rect 515 784 537 818
rect 537 784 549 818
rect 587 784 605 818
rect 605 784 621 818
rect 659 784 673 818
rect 673 784 693 818
rect 731 784 741 818
rect 741 784 765 818
rect 803 784 809 818
rect 809 784 837 818
rect 875 784 877 818
rect 877 784 909 818
rect 947 784 979 818
rect 979 784 981 818
rect 1019 784 1047 818
rect 1047 784 1053 818
rect 1091 784 1115 818
rect 1115 784 1125 818
rect 1163 784 1183 818
rect 1183 784 1197 818
rect 1235 784 1251 818
rect 1251 784 1269 818
rect 1307 784 1319 818
rect 1319 784 1341 818
rect 1379 784 1387 818
rect 1387 784 1413 818
rect 1451 784 1455 818
rect 1455 784 1485 818
rect 1523 784 1557 818
rect 1595 784 1625 818
rect 1625 784 1629 818
rect 1667 784 1693 818
rect 1693 784 1701 818
rect 1739 784 1761 818
rect 1761 784 1773 818
rect 1811 784 1829 818
rect 1829 784 1845 818
rect 1883 784 1897 818
rect 1897 784 1917 818
rect 1955 784 1965 818
rect 1965 784 1989 818
rect 2027 784 2033 818
rect 2033 784 2061 818
rect 2099 784 2101 818
rect 2101 784 2133 818
rect 2171 784 2203 818
rect 2203 784 2205 818
rect 2243 784 2271 818
rect 2271 784 2277 818
rect 2315 784 2339 818
rect 2339 784 2349 818
rect 2387 784 2407 818
rect 2407 784 2421 818
rect 2459 784 2475 818
rect 2475 784 2493 818
rect 2531 784 2543 818
rect 2543 784 2565 818
rect 2603 784 2611 818
rect 2611 784 2637 818
rect 2675 784 2679 818
rect 2679 784 2709 818
rect 2747 784 2781 818
rect 2819 784 2849 818
rect 2849 784 2853 818
rect 2891 784 2917 818
rect 2917 784 2925 818
rect 2963 784 2985 818
rect 2985 784 2997 818
rect 3035 784 3053 818
rect 3053 784 3069 818
rect 3233 784 3245 818
rect 3245 784 3267 818
rect 3305 784 3313 818
rect 3313 784 3339 818
rect 3377 784 3381 818
rect 3381 784 3411 818
rect 3449 784 3483 818
rect 3521 784 3551 818
rect 3551 784 3555 818
rect 3593 784 3619 818
rect 3619 784 3627 818
rect 3665 784 3687 818
rect 3687 784 3699 818
rect 3737 784 3755 818
rect 3755 784 3771 818
rect 3809 784 3823 818
rect 3823 784 3843 818
rect 3881 784 3891 818
rect 3891 784 3915 818
rect 3953 784 3959 818
rect 3959 784 3987 818
rect 4025 784 4027 818
rect 4027 784 4059 818
rect 4097 784 4129 818
rect 4129 784 4131 818
rect 4169 784 4197 818
rect 4197 784 4203 818
rect 4241 784 4265 818
rect 4265 784 4275 818
rect 4313 784 4333 818
rect 4333 784 4347 818
rect 4385 784 4401 818
rect 4401 784 4419 818
rect 4457 784 4469 818
rect 4469 784 4491 818
rect 4529 784 4537 818
rect 4537 784 4563 818
rect 4601 784 4605 818
rect 4605 784 4635 818
rect 4673 784 4707 818
rect 4745 784 4775 818
rect 4775 784 4779 818
rect 4817 784 4843 818
rect 4843 784 4851 818
rect 4889 784 4911 818
rect 4911 784 4923 818
rect 4961 784 4979 818
rect 4979 784 4995 818
rect 5033 784 5047 818
rect 5047 784 5067 818
rect 5105 784 5115 818
rect 5115 784 5139 818
rect 5177 784 5183 818
rect 5183 784 5211 818
rect 5249 784 5251 818
rect 5251 784 5283 818
rect 5321 784 5353 818
rect 5353 784 5355 818
rect 5393 784 5421 818
rect 5421 784 5427 818
rect 5465 784 5489 818
rect 5489 784 5499 818
rect 5537 784 5557 818
rect 5557 784 5571 818
rect 5609 784 5625 818
rect 5625 784 5643 818
rect 5681 784 5693 818
rect 5693 784 5715 818
rect 5753 784 5761 818
rect 5761 784 5787 818
rect 5825 784 5829 818
rect 5829 784 5859 818
rect 5897 784 5931 818
rect 5969 784 5999 818
rect 5999 784 6003 818
rect 6041 784 6067 818
rect 6067 784 6075 818
rect 6113 784 6135 818
rect 6135 784 6147 818
rect 6185 784 6203 818
rect 6203 784 6219 818
rect 9388 837 9422 871
rect 6273 768 6307 801
rect 6273 767 6307 768
rect 9460 837 9494 871
rect 12538 837 12572 871
rect 3088 707 3122 741
rect 3160 707 3194 741
rect 6383 758 6395 792
rect 6395 758 6417 792
rect 6455 758 6463 792
rect 6463 758 6489 792
rect 6527 758 6531 792
rect 6531 758 6561 792
rect 6599 758 6633 792
rect 6671 758 6701 792
rect 6701 758 6705 792
rect 6743 758 6769 792
rect 6769 758 6777 792
rect 6815 758 6837 792
rect 6837 758 6849 792
rect 6887 758 6905 792
rect 6905 758 6921 792
rect 6959 758 6973 792
rect 6973 758 6993 792
rect 7031 758 7041 792
rect 7041 758 7065 792
rect 7103 758 7109 792
rect 7109 758 7137 792
rect 7175 758 7177 792
rect 7177 758 7209 792
rect 7247 758 7279 792
rect 7279 758 7281 792
rect 7319 758 7347 792
rect 7347 758 7353 792
rect 7391 758 7415 792
rect 7415 758 7425 792
rect 7463 758 7483 792
rect 7483 758 7497 792
rect 7535 758 7551 792
rect 7551 758 7569 792
rect 7607 758 7619 792
rect 7619 758 7641 792
rect 7679 758 7687 792
rect 7687 758 7713 792
rect 7751 758 7755 792
rect 7755 758 7785 792
rect 7823 758 7857 792
rect 7895 758 7925 792
rect 7925 758 7929 792
rect 7967 758 7993 792
rect 7993 758 8001 792
rect 8039 758 8061 792
rect 8061 758 8073 792
rect 8111 758 8129 792
rect 8129 758 8145 792
rect 8183 758 8197 792
rect 8197 758 8217 792
rect 8255 758 8265 792
rect 8265 758 8289 792
rect 8327 758 8333 792
rect 8333 758 8361 792
rect 8399 758 8401 792
rect 8401 758 8433 792
rect 8471 758 8503 792
rect 8503 758 8505 792
rect 8543 758 8571 792
rect 8571 758 8577 792
rect 8615 758 8639 792
rect 8639 758 8649 792
rect 8687 758 8707 792
rect 8707 758 8721 792
rect 8759 758 8775 792
rect 8775 758 8793 792
rect 8831 758 8843 792
rect 8843 758 8865 792
rect 8903 758 8911 792
rect 8911 758 8937 792
rect 8975 758 8979 792
rect 8979 758 9009 792
rect 9047 758 9081 792
rect 9119 758 9149 792
rect 9149 758 9153 792
rect 9191 758 9217 792
rect 9217 758 9225 792
rect 9263 758 9285 792
rect 9285 758 9297 792
rect 9335 758 9353 792
rect 9353 758 9369 792
rect 12610 837 12644 871
rect 15688 837 15722 871
rect 6273 723 6307 725
rect 6273 691 6307 723
rect 9533 758 9545 792
rect 9545 758 9567 792
rect 9605 758 9613 792
rect 9613 758 9639 792
rect 9677 758 9681 792
rect 9681 758 9711 792
rect 9749 758 9783 792
rect 9821 758 9851 792
rect 9851 758 9855 792
rect 9893 758 9919 792
rect 9919 758 9927 792
rect 9965 758 9987 792
rect 9987 758 9999 792
rect 10037 758 10055 792
rect 10055 758 10071 792
rect 10109 758 10123 792
rect 10123 758 10143 792
rect 10181 758 10191 792
rect 10191 758 10215 792
rect 10253 758 10259 792
rect 10259 758 10287 792
rect 10325 758 10327 792
rect 10327 758 10359 792
rect 10397 758 10429 792
rect 10429 758 10431 792
rect 10469 758 10497 792
rect 10497 758 10503 792
rect 10541 758 10565 792
rect 10565 758 10575 792
rect 10613 758 10633 792
rect 10633 758 10647 792
rect 10685 758 10701 792
rect 10701 758 10719 792
rect 10757 758 10769 792
rect 10769 758 10791 792
rect 10829 758 10837 792
rect 10837 758 10863 792
rect 10901 758 10905 792
rect 10905 758 10935 792
rect 10973 758 11007 792
rect 11045 758 11075 792
rect 11075 758 11079 792
rect 11117 758 11143 792
rect 11143 758 11151 792
rect 11189 758 11211 792
rect 11211 758 11223 792
rect 11261 758 11279 792
rect 11279 758 11295 792
rect 11333 758 11347 792
rect 11347 758 11367 792
rect 11405 758 11415 792
rect 11415 758 11439 792
rect 11477 758 11483 792
rect 11483 758 11511 792
rect 11549 758 11551 792
rect 11551 758 11583 792
rect 11621 758 11653 792
rect 11653 758 11655 792
rect 11693 758 11721 792
rect 11721 758 11727 792
rect 11765 758 11789 792
rect 11789 758 11799 792
rect 11837 758 11857 792
rect 11857 758 11871 792
rect 11909 758 11925 792
rect 11925 758 11943 792
rect 11981 758 11993 792
rect 11993 758 12015 792
rect 12053 758 12061 792
rect 12061 758 12087 792
rect 12125 758 12129 792
rect 12129 758 12159 792
rect 12197 758 12231 792
rect 12269 758 12299 792
rect 12299 758 12303 792
rect 12341 758 12367 792
rect 12367 758 12375 792
rect 12413 758 12435 792
rect 12435 758 12447 792
rect 12485 758 12503 792
rect 12503 758 12519 792
rect 15760 837 15794 871
rect 18838 837 18872 871
rect 12683 758 12695 792
rect 12695 758 12717 792
rect 12755 758 12763 792
rect 12763 758 12789 792
rect 12827 758 12831 792
rect 12831 758 12861 792
rect 12899 758 12933 792
rect 12971 758 13001 792
rect 13001 758 13005 792
rect 13043 758 13069 792
rect 13069 758 13077 792
rect 13115 758 13137 792
rect 13137 758 13149 792
rect 13187 758 13205 792
rect 13205 758 13221 792
rect 13259 758 13273 792
rect 13273 758 13293 792
rect 13331 758 13341 792
rect 13341 758 13365 792
rect 13403 758 13409 792
rect 13409 758 13437 792
rect 13475 758 13477 792
rect 13477 758 13509 792
rect 13547 758 13579 792
rect 13579 758 13581 792
rect 13619 758 13647 792
rect 13647 758 13653 792
rect 13691 758 13715 792
rect 13715 758 13725 792
rect 13763 758 13783 792
rect 13783 758 13797 792
rect 13835 758 13851 792
rect 13851 758 13869 792
rect 13907 758 13919 792
rect 13919 758 13941 792
rect 13979 758 13987 792
rect 13987 758 14013 792
rect 14051 758 14055 792
rect 14055 758 14085 792
rect 14123 758 14157 792
rect 14195 758 14225 792
rect 14225 758 14229 792
rect 14267 758 14293 792
rect 14293 758 14301 792
rect 14339 758 14361 792
rect 14361 758 14373 792
rect 14411 758 14429 792
rect 14429 758 14445 792
rect 14483 758 14497 792
rect 14497 758 14517 792
rect 14555 758 14565 792
rect 14565 758 14589 792
rect 14627 758 14633 792
rect 14633 758 14661 792
rect 14699 758 14701 792
rect 14701 758 14733 792
rect 14771 758 14803 792
rect 14803 758 14805 792
rect 14843 758 14871 792
rect 14871 758 14877 792
rect 14915 758 14939 792
rect 14939 758 14949 792
rect 14987 758 15007 792
rect 15007 758 15021 792
rect 15059 758 15075 792
rect 15075 758 15093 792
rect 15131 758 15143 792
rect 15143 758 15165 792
rect 15203 758 15211 792
rect 15211 758 15237 792
rect 15275 758 15279 792
rect 15279 758 15309 792
rect 15347 758 15381 792
rect 15419 758 15449 792
rect 15449 758 15453 792
rect 15491 758 15517 792
rect 15517 758 15525 792
rect 15563 758 15585 792
rect 15585 758 15597 792
rect 15635 758 15653 792
rect 15653 758 15669 792
rect 18910 837 18944 871
rect 21988 837 22022 871
rect 15833 758 15845 792
rect 15845 758 15867 792
rect 15905 758 15913 792
rect 15913 758 15939 792
rect 15977 758 15981 792
rect 15981 758 16011 792
rect 16049 758 16083 792
rect 16121 758 16151 792
rect 16151 758 16155 792
rect 16193 758 16219 792
rect 16219 758 16227 792
rect 16265 758 16287 792
rect 16287 758 16299 792
rect 16337 758 16355 792
rect 16355 758 16371 792
rect 16409 758 16423 792
rect 16423 758 16443 792
rect 16481 758 16491 792
rect 16491 758 16515 792
rect 16553 758 16559 792
rect 16559 758 16587 792
rect 16625 758 16627 792
rect 16627 758 16659 792
rect 16697 758 16729 792
rect 16729 758 16731 792
rect 16769 758 16797 792
rect 16797 758 16803 792
rect 16841 758 16865 792
rect 16865 758 16875 792
rect 16913 758 16933 792
rect 16933 758 16947 792
rect 16985 758 17001 792
rect 17001 758 17019 792
rect 17057 758 17069 792
rect 17069 758 17091 792
rect 17129 758 17137 792
rect 17137 758 17163 792
rect 17201 758 17205 792
rect 17205 758 17235 792
rect 17273 758 17307 792
rect 17345 758 17375 792
rect 17375 758 17379 792
rect 17417 758 17443 792
rect 17443 758 17451 792
rect 17489 758 17511 792
rect 17511 758 17523 792
rect 17561 758 17579 792
rect 17579 758 17595 792
rect 17633 758 17647 792
rect 17647 758 17667 792
rect 17705 758 17715 792
rect 17715 758 17739 792
rect 17777 758 17783 792
rect 17783 758 17811 792
rect 17849 758 17851 792
rect 17851 758 17883 792
rect 17921 758 17953 792
rect 17953 758 17955 792
rect 17993 758 18021 792
rect 18021 758 18027 792
rect 18065 758 18089 792
rect 18089 758 18099 792
rect 18137 758 18157 792
rect 18157 758 18171 792
rect 18209 758 18225 792
rect 18225 758 18243 792
rect 18281 758 18293 792
rect 18293 758 18315 792
rect 18353 758 18361 792
rect 18361 758 18387 792
rect 18425 758 18429 792
rect 18429 758 18459 792
rect 18497 758 18531 792
rect 18569 758 18599 792
rect 18599 758 18603 792
rect 18641 758 18667 792
rect 18667 758 18675 792
rect 18713 758 18735 792
rect 18735 758 18747 792
rect 18785 758 18803 792
rect 18803 758 18819 792
rect 22060 837 22094 871
rect 18983 758 18995 792
rect 18995 758 19017 792
rect 19055 758 19063 792
rect 19063 758 19089 792
rect 19127 758 19131 792
rect 19131 758 19161 792
rect 19199 758 19233 792
rect 19271 758 19301 792
rect 19301 758 19305 792
rect 19343 758 19369 792
rect 19369 758 19377 792
rect 19415 758 19437 792
rect 19437 758 19449 792
rect 19487 758 19505 792
rect 19505 758 19521 792
rect 19559 758 19573 792
rect 19573 758 19593 792
rect 19631 758 19641 792
rect 19641 758 19665 792
rect 19703 758 19709 792
rect 19709 758 19737 792
rect 19775 758 19777 792
rect 19777 758 19809 792
rect 19847 758 19879 792
rect 19879 758 19881 792
rect 19919 758 19947 792
rect 19947 758 19953 792
rect 19991 758 20015 792
rect 20015 758 20025 792
rect 20063 758 20083 792
rect 20083 758 20097 792
rect 20135 758 20151 792
rect 20151 758 20169 792
rect 20207 758 20219 792
rect 20219 758 20241 792
rect 20279 758 20287 792
rect 20287 758 20313 792
rect 20351 758 20355 792
rect 20355 758 20385 792
rect 20423 758 20457 792
rect 20495 758 20525 792
rect 20525 758 20529 792
rect 20567 758 20593 792
rect 20593 758 20601 792
rect 20639 758 20661 792
rect 20661 758 20673 792
rect 20711 758 20729 792
rect 20729 758 20745 792
rect 20783 758 20797 792
rect 20797 758 20817 792
rect 20855 758 20865 792
rect 20865 758 20889 792
rect 20927 758 20933 792
rect 20933 758 20961 792
rect 20999 758 21001 792
rect 21001 758 21033 792
rect 21071 758 21103 792
rect 21103 758 21105 792
rect 21143 758 21171 792
rect 21171 758 21177 792
rect 21215 758 21239 792
rect 21239 758 21249 792
rect 21287 758 21307 792
rect 21307 758 21321 792
rect 21359 758 21375 792
rect 21375 758 21393 792
rect 21431 758 21443 792
rect 21443 758 21465 792
rect 21503 758 21511 792
rect 21511 758 21537 792
rect 21575 758 21579 792
rect 21579 758 21609 792
rect 21647 758 21681 792
rect 21719 758 21749 792
rect 21749 758 21753 792
rect 21791 758 21817 792
rect 21817 758 21825 792
rect 21863 758 21885 792
rect 21885 758 21897 792
rect 21935 758 21953 792
rect 21953 758 21969 792
rect 22248 835 22282 836
rect 22248 802 22282 835
rect 22366 824 22390 858
rect 22390 824 22400 858
rect 22438 824 22458 858
rect 22458 824 22472 858
rect 22510 824 22526 858
rect 22526 824 22544 858
rect 22582 824 22594 858
rect 22594 824 22616 858
rect 22654 824 22662 858
rect 22662 824 22688 858
rect 22726 824 22730 858
rect 22730 824 22760 858
rect 22798 824 22832 858
rect 22870 824 22900 858
rect 22900 824 22904 858
rect 22942 824 22968 858
rect 22968 824 22976 858
rect 23014 824 23036 858
rect 23036 824 23048 858
rect 23086 824 23104 858
rect 23104 824 23120 858
rect 23158 824 23172 858
rect 23172 824 23192 858
rect 23230 824 23240 858
rect 23240 824 23264 858
rect 23302 824 23308 858
rect 23308 824 23336 858
rect 23374 824 23376 858
rect 23376 824 23408 858
rect 23446 824 23478 858
rect 23478 824 23480 858
rect 23518 824 23546 858
rect 23546 824 23552 858
rect 23590 824 23614 858
rect 23614 824 23624 858
rect 23662 824 23682 858
rect 23682 824 23696 858
rect 23734 824 23750 858
rect 23750 824 23768 858
rect 23806 824 23818 858
rect 23818 824 23840 858
rect 23878 824 23886 858
rect 23886 824 23912 858
rect 23950 824 23954 858
rect 23954 824 23984 858
rect 24022 824 24056 858
rect 24094 824 24124 858
rect 24124 824 24128 858
rect 24166 824 24192 858
rect 24192 824 24200 858
rect 24238 824 24260 858
rect 24260 824 24272 858
rect 24310 824 24328 858
rect 24328 824 24344 858
rect 22248 729 22282 760
rect 22248 726 22282 729
rect 83 628 95 662
rect 95 628 117 662
rect 155 628 163 662
rect 163 628 189 662
rect 227 628 231 662
rect 231 628 261 662
rect 299 628 333 662
rect 371 628 401 662
rect 401 628 405 662
rect 443 628 469 662
rect 469 628 477 662
rect 515 628 537 662
rect 537 628 549 662
rect 587 628 605 662
rect 605 628 621 662
rect 659 628 673 662
rect 673 628 693 662
rect 731 628 741 662
rect 741 628 765 662
rect 803 628 809 662
rect 809 628 837 662
rect 875 628 877 662
rect 877 628 909 662
rect 947 628 979 662
rect 979 628 981 662
rect 1019 628 1047 662
rect 1047 628 1053 662
rect 1091 628 1115 662
rect 1115 628 1125 662
rect 1163 628 1183 662
rect 1183 628 1197 662
rect 1235 628 1251 662
rect 1251 628 1269 662
rect 1307 628 1319 662
rect 1319 628 1341 662
rect 1379 628 1387 662
rect 1387 628 1413 662
rect 1451 628 1455 662
rect 1455 628 1485 662
rect 1523 628 1557 662
rect 1595 628 1625 662
rect 1625 628 1629 662
rect 1667 628 1693 662
rect 1693 628 1701 662
rect 1739 628 1761 662
rect 1761 628 1773 662
rect 1811 628 1829 662
rect 1829 628 1845 662
rect 1883 628 1897 662
rect 1897 628 1917 662
rect 1955 628 1965 662
rect 1965 628 1989 662
rect 2027 628 2033 662
rect 2033 628 2061 662
rect 2099 628 2101 662
rect 2101 628 2133 662
rect 2171 628 2203 662
rect 2203 628 2205 662
rect 2243 628 2271 662
rect 2271 628 2277 662
rect 2315 628 2339 662
rect 2339 628 2349 662
rect 2387 628 2407 662
rect 2407 628 2421 662
rect 2459 628 2475 662
rect 2475 628 2493 662
rect 2531 628 2543 662
rect 2543 628 2565 662
rect 2603 628 2611 662
rect 2611 628 2637 662
rect 2675 628 2679 662
rect 2679 628 2709 662
rect 2747 628 2781 662
rect 2819 628 2849 662
rect 2849 628 2853 662
rect 2891 628 2917 662
rect 2917 628 2925 662
rect 2963 628 2985 662
rect 2985 628 2997 662
rect 3035 628 3053 662
rect 3053 628 3069 662
rect 3233 628 3245 662
rect 3245 628 3267 662
rect 3305 628 3313 662
rect 3313 628 3339 662
rect 3377 628 3381 662
rect 3381 628 3411 662
rect 3449 628 3483 662
rect 3521 628 3551 662
rect 3551 628 3555 662
rect 3593 628 3619 662
rect 3619 628 3627 662
rect 3665 628 3687 662
rect 3687 628 3699 662
rect 3737 628 3755 662
rect 3755 628 3771 662
rect 3809 628 3823 662
rect 3823 628 3843 662
rect 3881 628 3891 662
rect 3891 628 3915 662
rect 3953 628 3959 662
rect 3959 628 3987 662
rect 4025 628 4027 662
rect 4027 628 4059 662
rect 4097 628 4129 662
rect 4129 628 4131 662
rect 4169 628 4197 662
rect 4197 628 4203 662
rect 4241 628 4265 662
rect 4265 628 4275 662
rect 4313 628 4333 662
rect 4333 628 4347 662
rect 4385 628 4401 662
rect 4401 628 4419 662
rect 4457 628 4469 662
rect 4469 628 4491 662
rect 4529 628 4537 662
rect 4537 628 4563 662
rect 4601 628 4605 662
rect 4605 628 4635 662
rect 4673 628 4707 662
rect 4745 628 4775 662
rect 4775 628 4779 662
rect 4817 628 4843 662
rect 4843 628 4851 662
rect 4889 628 4911 662
rect 4911 628 4923 662
rect 4961 628 4979 662
rect 4979 628 4995 662
rect 5033 628 5047 662
rect 5047 628 5067 662
rect 5105 628 5115 662
rect 5115 628 5139 662
rect 5177 628 5183 662
rect 5183 628 5211 662
rect 5249 628 5251 662
rect 5251 628 5283 662
rect 5321 628 5353 662
rect 5353 628 5355 662
rect 5393 628 5421 662
rect 5421 628 5427 662
rect 5465 628 5489 662
rect 5489 628 5499 662
rect 5537 628 5557 662
rect 5557 628 5571 662
rect 5609 628 5625 662
rect 5625 628 5643 662
rect 5681 628 5693 662
rect 5693 628 5715 662
rect 5753 628 5761 662
rect 5761 628 5787 662
rect 5825 628 5829 662
rect 5829 628 5859 662
rect 5897 628 5931 662
rect 5969 628 5999 662
rect 5999 628 6003 662
rect 6041 628 6067 662
rect 6067 628 6075 662
rect 6113 628 6135 662
rect 6135 628 6147 662
rect 6185 628 6203 662
rect 6203 628 6219 662
rect 9388 681 9422 715
rect 9460 681 9494 715
rect 12538 681 12572 715
rect 12610 681 12644 715
rect 15688 681 15722 715
rect 15760 681 15794 715
rect 18838 681 18872 715
rect 18910 681 18944 715
rect 21988 681 22022 715
rect 22060 681 22094 715
rect 22366 668 22390 702
rect 22390 668 22400 702
rect 22438 668 22458 702
rect 22458 668 22472 702
rect 22510 668 22526 702
rect 22526 668 22544 702
rect 22582 668 22594 702
rect 22594 668 22616 702
rect 22654 668 22662 702
rect 22662 668 22688 702
rect 22726 668 22730 702
rect 22730 668 22760 702
rect 22798 668 22832 702
rect 22870 668 22900 702
rect 22900 668 22904 702
rect 22942 668 22968 702
rect 22968 668 22976 702
rect 23014 668 23036 702
rect 23036 668 23048 702
rect 23086 668 23104 702
rect 23104 668 23120 702
rect 23158 668 23172 702
rect 23172 668 23192 702
rect 23230 668 23240 702
rect 23240 668 23264 702
rect 23302 668 23308 702
rect 23308 668 23336 702
rect 23374 668 23376 702
rect 23376 668 23408 702
rect 23446 668 23478 702
rect 23478 668 23480 702
rect 23518 668 23546 702
rect 23546 668 23552 702
rect 23590 668 23614 702
rect 23614 668 23624 702
rect 23662 668 23682 702
rect 23682 668 23696 702
rect 23734 668 23750 702
rect 23750 668 23768 702
rect 23806 668 23818 702
rect 23818 668 23840 702
rect 23878 668 23886 702
rect 23886 668 23912 702
rect 23950 668 23954 702
rect 23954 668 23984 702
rect 24022 668 24056 702
rect 24094 668 24124 702
rect 24124 668 24128 702
rect 24166 668 24192 702
rect 24192 668 24200 702
rect 24238 668 24260 702
rect 24260 668 24272 702
rect 24310 668 24328 702
rect 24328 668 24344 702
rect 6383 602 6395 636
rect 6395 602 6417 636
rect 6455 602 6463 636
rect 6463 602 6489 636
rect 6527 602 6531 636
rect 6531 602 6561 636
rect 6599 602 6633 636
rect 6671 602 6701 636
rect 6701 602 6705 636
rect 6743 602 6769 636
rect 6769 602 6777 636
rect 6815 602 6837 636
rect 6837 602 6849 636
rect 6887 602 6905 636
rect 6905 602 6921 636
rect 6959 602 6973 636
rect 6973 602 6993 636
rect 7031 602 7041 636
rect 7041 602 7065 636
rect 7103 602 7109 636
rect 7109 602 7137 636
rect 7175 602 7177 636
rect 7177 602 7209 636
rect 7247 602 7279 636
rect 7279 602 7281 636
rect 7319 602 7347 636
rect 7347 602 7353 636
rect 7391 602 7415 636
rect 7415 602 7425 636
rect 7463 602 7483 636
rect 7483 602 7497 636
rect 7535 602 7551 636
rect 7551 602 7569 636
rect 7607 602 7619 636
rect 7619 602 7641 636
rect 7679 602 7687 636
rect 7687 602 7713 636
rect 7751 602 7755 636
rect 7755 602 7785 636
rect 7823 602 7857 636
rect 7895 602 7925 636
rect 7925 602 7929 636
rect 7967 602 7993 636
rect 7993 602 8001 636
rect 8039 602 8061 636
rect 8061 602 8073 636
rect 8111 602 8129 636
rect 8129 602 8145 636
rect 8183 602 8197 636
rect 8197 602 8217 636
rect 8255 602 8265 636
rect 8265 602 8289 636
rect 8327 602 8333 636
rect 8333 602 8361 636
rect 8399 602 8401 636
rect 8401 602 8433 636
rect 8471 602 8503 636
rect 8503 602 8505 636
rect 8543 602 8571 636
rect 8571 602 8577 636
rect 8615 602 8639 636
rect 8639 602 8649 636
rect 8687 602 8707 636
rect 8707 602 8721 636
rect 8759 602 8775 636
rect 8775 602 8793 636
rect 8831 602 8843 636
rect 8843 602 8865 636
rect 8903 602 8911 636
rect 8911 602 8937 636
rect 8975 602 8979 636
rect 8979 602 9009 636
rect 9047 602 9081 636
rect 9119 602 9149 636
rect 9149 602 9153 636
rect 9191 602 9217 636
rect 9217 602 9225 636
rect 9263 602 9285 636
rect 9285 602 9297 636
rect 9335 602 9353 636
rect 9353 602 9369 636
rect 9533 602 9545 636
rect 9545 602 9567 636
rect 9605 602 9613 636
rect 9613 602 9639 636
rect 9677 602 9681 636
rect 9681 602 9711 636
rect 9749 602 9783 636
rect 9821 602 9851 636
rect 9851 602 9855 636
rect 9893 602 9919 636
rect 9919 602 9927 636
rect 9965 602 9987 636
rect 9987 602 9999 636
rect 10037 602 10055 636
rect 10055 602 10071 636
rect 10109 602 10123 636
rect 10123 602 10143 636
rect 10181 602 10191 636
rect 10191 602 10215 636
rect 10253 602 10259 636
rect 10259 602 10287 636
rect 10325 602 10327 636
rect 10327 602 10359 636
rect 10397 602 10429 636
rect 10429 602 10431 636
rect 10469 602 10497 636
rect 10497 602 10503 636
rect 10541 602 10565 636
rect 10565 602 10575 636
rect 10613 602 10633 636
rect 10633 602 10647 636
rect 10685 602 10701 636
rect 10701 602 10719 636
rect 10757 602 10769 636
rect 10769 602 10791 636
rect 10829 602 10837 636
rect 10837 602 10863 636
rect 10901 602 10905 636
rect 10905 602 10935 636
rect 10973 602 11007 636
rect 11045 602 11075 636
rect 11075 602 11079 636
rect 11117 602 11143 636
rect 11143 602 11151 636
rect 11189 602 11211 636
rect 11211 602 11223 636
rect 11261 602 11279 636
rect 11279 602 11295 636
rect 11333 602 11347 636
rect 11347 602 11367 636
rect 11405 602 11415 636
rect 11415 602 11439 636
rect 11477 602 11483 636
rect 11483 602 11511 636
rect 11549 602 11551 636
rect 11551 602 11583 636
rect 11621 602 11653 636
rect 11653 602 11655 636
rect 11693 602 11721 636
rect 11721 602 11727 636
rect 11765 602 11789 636
rect 11789 602 11799 636
rect 11837 602 11857 636
rect 11857 602 11871 636
rect 11909 602 11925 636
rect 11925 602 11943 636
rect 11981 602 11993 636
rect 11993 602 12015 636
rect 12053 602 12061 636
rect 12061 602 12087 636
rect 12125 602 12129 636
rect 12129 602 12159 636
rect 12197 602 12231 636
rect 12269 602 12299 636
rect 12299 602 12303 636
rect 12341 602 12367 636
rect 12367 602 12375 636
rect 12413 602 12435 636
rect 12435 602 12447 636
rect 12485 602 12503 636
rect 12503 602 12519 636
rect 12683 602 12695 636
rect 12695 602 12717 636
rect 12755 602 12763 636
rect 12763 602 12789 636
rect 12827 602 12831 636
rect 12831 602 12861 636
rect 12899 602 12933 636
rect 12971 602 13001 636
rect 13001 602 13005 636
rect 13043 602 13069 636
rect 13069 602 13077 636
rect 13115 602 13137 636
rect 13137 602 13149 636
rect 13187 602 13205 636
rect 13205 602 13221 636
rect 13259 602 13273 636
rect 13273 602 13293 636
rect 13331 602 13341 636
rect 13341 602 13365 636
rect 13403 602 13409 636
rect 13409 602 13437 636
rect 13475 602 13477 636
rect 13477 602 13509 636
rect 13547 602 13579 636
rect 13579 602 13581 636
rect 13619 602 13647 636
rect 13647 602 13653 636
rect 13691 602 13715 636
rect 13715 602 13725 636
rect 13763 602 13783 636
rect 13783 602 13797 636
rect 13835 602 13851 636
rect 13851 602 13869 636
rect 13907 602 13919 636
rect 13919 602 13941 636
rect 13979 602 13987 636
rect 13987 602 14013 636
rect 14051 602 14055 636
rect 14055 602 14085 636
rect 14123 602 14157 636
rect 14195 602 14225 636
rect 14225 602 14229 636
rect 14267 602 14293 636
rect 14293 602 14301 636
rect 14339 602 14361 636
rect 14361 602 14373 636
rect 14411 602 14429 636
rect 14429 602 14445 636
rect 14483 602 14497 636
rect 14497 602 14517 636
rect 14555 602 14565 636
rect 14565 602 14589 636
rect 14627 602 14633 636
rect 14633 602 14661 636
rect 14699 602 14701 636
rect 14701 602 14733 636
rect 14771 602 14803 636
rect 14803 602 14805 636
rect 14843 602 14871 636
rect 14871 602 14877 636
rect 14915 602 14939 636
rect 14939 602 14949 636
rect 14987 602 15007 636
rect 15007 602 15021 636
rect 15059 602 15075 636
rect 15075 602 15093 636
rect 15131 602 15143 636
rect 15143 602 15165 636
rect 15203 602 15211 636
rect 15211 602 15237 636
rect 15275 602 15279 636
rect 15279 602 15309 636
rect 15347 602 15381 636
rect 15419 602 15449 636
rect 15449 602 15453 636
rect 15491 602 15517 636
rect 15517 602 15525 636
rect 15563 602 15585 636
rect 15585 602 15597 636
rect 15635 602 15653 636
rect 15653 602 15669 636
rect 15833 602 15845 636
rect 15845 602 15867 636
rect 15905 602 15913 636
rect 15913 602 15939 636
rect 15977 602 15981 636
rect 15981 602 16011 636
rect 16049 602 16083 636
rect 16121 602 16151 636
rect 16151 602 16155 636
rect 16193 602 16219 636
rect 16219 602 16227 636
rect 16265 602 16287 636
rect 16287 602 16299 636
rect 16337 602 16355 636
rect 16355 602 16371 636
rect 16409 602 16423 636
rect 16423 602 16443 636
rect 16481 602 16491 636
rect 16491 602 16515 636
rect 16553 602 16559 636
rect 16559 602 16587 636
rect 16625 602 16627 636
rect 16627 602 16659 636
rect 16697 602 16729 636
rect 16729 602 16731 636
rect 16769 602 16797 636
rect 16797 602 16803 636
rect 16841 602 16865 636
rect 16865 602 16875 636
rect 16913 602 16933 636
rect 16933 602 16947 636
rect 16985 602 17001 636
rect 17001 602 17019 636
rect 17057 602 17069 636
rect 17069 602 17091 636
rect 17129 602 17137 636
rect 17137 602 17163 636
rect 17201 602 17205 636
rect 17205 602 17235 636
rect 17273 602 17307 636
rect 17345 602 17375 636
rect 17375 602 17379 636
rect 17417 602 17443 636
rect 17443 602 17451 636
rect 17489 602 17511 636
rect 17511 602 17523 636
rect 17561 602 17579 636
rect 17579 602 17595 636
rect 17633 602 17647 636
rect 17647 602 17667 636
rect 17705 602 17715 636
rect 17715 602 17739 636
rect 17777 602 17783 636
rect 17783 602 17811 636
rect 17849 602 17851 636
rect 17851 602 17883 636
rect 17921 602 17953 636
rect 17953 602 17955 636
rect 17993 602 18021 636
rect 18021 602 18027 636
rect 18065 602 18089 636
rect 18089 602 18099 636
rect 18137 602 18157 636
rect 18157 602 18171 636
rect 18209 602 18225 636
rect 18225 602 18243 636
rect 18281 602 18293 636
rect 18293 602 18315 636
rect 18353 602 18361 636
rect 18361 602 18387 636
rect 18425 602 18429 636
rect 18429 602 18459 636
rect 18497 602 18531 636
rect 18569 602 18599 636
rect 18599 602 18603 636
rect 18641 602 18667 636
rect 18667 602 18675 636
rect 18713 602 18735 636
rect 18735 602 18747 636
rect 18785 602 18803 636
rect 18803 602 18819 636
rect 18983 602 18995 636
rect 18995 602 19017 636
rect 19055 602 19063 636
rect 19063 602 19089 636
rect 19127 602 19131 636
rect 19131 602 19161 636
rect 19199 602 19233 636
rect 19271 602 19301 636
rect 19301 602 19305 636
rect 19343 602 19369 636
rect 19369 602 19377 636
rect 19415 602 19437 636
rect 19437 602 19449 636
rect 19487 602 19505 636
rect 19505 602 19521 636
rect 19559 602 19573 636
rect 19573 602 19593 636
rect 19631 602 19641 636
rect 19641 602 19665 636
rect 19703 602 19709 636
rect 19709 602 19737 636
rect 19775 602 19777 636
rect 19777 602 19809 636
rect 19847 602 19879 636
rect 19879 602 19881 636
rect 19919 602 19947 636
rect 19947 602 19953 636
rect 19991 602 20015 636
rect 20015 602 20025 636
rect 20063 602 20083 636
rect 20083 602 20097 636
rect 20135 602 20151 636
rect 20151 602 20169 636
rect 20207 602 20219 636
rect 20219 602 20241 636
rect 20279 602 20287 636
rect 20287 602 20313 636
rect 20351 602 20355 636
rect 20355 602 20385 636
rect 20423 602 20457 636
rect 20495 602 20525 636
rect 20525 602 20529 636
rect 20567 602 20593 636
rect 20593 602 20601 636
rect 20639 602 20661 636
rect 20661 602 20673 636
rect 20711 602 20729 636
rect 20729 602 20745 636
rect 20783 602 20797 636
rect 20797 602 20817 636
rect 20855 602 20865 636
rect 20865 602 20889 636
rect 20927 602 20933 636
rect 20933 602 20961 636
rect 20999 602 21001 636
rect 21001 602 21033 636
rect 21071 602 21103 636
rect 21103 602 21105 636
rect 21143 602 21171 636
rect 21171 602 21177 636
rect 21215 602 21239 636
rect 21239 602 21249 636
rect 21287 602 21307 636
rect 21307 602 21321 636
rect 21359 602 21375 636
rect 21375 602 21393 636
rect 21431 602 21443 636
rect 21443 602 21465 636
rect 21503 602 21511 636
rect 21511 602 21537 636
rect 21575 602 21579 636
rect 21579 602 21609 636
rect 21647 602 21681 636
rect 21719 602 21749 636
rect 21749 602 21753 636
rect 21791 602 21817 636
rect 21817 602 21825 636
rect 21863 602 21885 636
rect 21885 602 21897 636
rect 21935 602 21953 636
rect 21953 602 21969 636
<< metal1 >>
tri 22426 2112 22429 2115 se
rect 22429 2112 22436 2115
rect 22354 2106 22436 2112
rect 22354 2072 22366 2106
rect 22400 2072 22436 2106
rect 22354 2066 22436 2072
tri 22426 2063 22429 2066 ne
rect 22429 2063 22436 2066
rect 22488 2063 22504 2115
rect 22556 2063 22572 2115
rect 22624 2063 22640 2115
rect 22692 2063 22708 2115
rect 22760 2063 22776 2115
rect 22828 2106 22844 2115
rect 22896 2106 22912 2115
rect 22964 2106 22980 2115
rect 23032 2106 23048 2115
rect 23100 2106 23116 2115
rect 23168 2106 23183 2115
rect 23235 2106 23250 2115
rect 23302 2112 23308 2115
tri 23308 2112 23311 2115 sw
rect 23302 2106 24356 2112
rect 22832 2072 22844 2106
rect 22904 2072 22912 2106
rect 22976 2072 22980 2106
rect 23336 2072 23374 2106
rect 23408 2072 23446 2106
rect 23480 2072 23518 2106
rect 23552 2072 23590 2106
rect 23624 2072 23662 2106
rect 23696 2072 23734 2106
rect 23768 2072 23806 2106
rect 23840 2072 23878 2106
rect 23912 2072 23950 2106
rect 23984 2072 24022 2106
rect 24056 2072 24094 2106
rect 24128 2072 24166 2106
rect 24200 2072 24238 2106
rect 24272 2072 24310 2106
rect 24344 2072 24356 2106
rect 22828 2063 22844 2072
rect 22896 2063 22912 2072
rect 22964 2063 22980 2072
rect 23032 2063 23048 2072
rect 23100 2063 23116 2072
rect 23168 2063 23183 2072
rect 23235 2063 23250 2072
rect 23302 2066 24356 2072
rect 23302 2063 23308 2066
tri 23308 2063 23311 2066 nw
rect 22236 2055 22288 2061
rect 22236 1991 22288 2003
tri 23398 1956 23401 1959 se
rect 23401 1956 23407 1959
rect 22236 1927 22288 1939
rect 22354 1950 23407 1956
rect 23459 1950 23478 1959
rect 23530 1950 23549 1959
rect 23601 1950 23620 1959
rect 23672 1950 23691 1959
rect 23743 1950 23762 1959
rect 23814 1950 23833 1959
rect 23885 1950 23904 1959
rect 23956 1950 23975 1959
rect 24027 1950 24046 1959
rect 24098 1956 24104 1959
tri 24104 1956 24107 1959 sw
rect 24098 1950 24356 1956
rect 22354 1916 22366 1950
rect 22400 1916 22438 1950
rect 22472 1916 22510 1950
rect 22544 1916 22582 1950
rect 22616 1916 22654 1950
rect 22688 1916 22726 1950
rect 22760 1916 22798 1950
rect 22832 1916 22870 1950
rect 22904 1916 22942 1950
rect 22976 1916 23014 1950
rect 23048 1916 23086 1950
rect 23120 1916 23158 1950
rect 23192 1916 23230 1950
rect 23264 1916 23302 1950
rect 23336 1916 23374 1950
rect 24128 1916 24166 1950
rect 24200 1916 24238 1950
rect 24272 1916 24310 1950
rect 24344 1916 24356 1950
rect 22354 1910 23407 1916
tri 23398 1907 23401 1910 ne
rect 23401 1907 23407 1910
rect 23459 1907 23478 1916
rect 23530 1907 23549 1916
rect 23601 1907 23620 1916
rect 23672 1907 23691 1916
rect 23743 1907 23762 1916
rect 23814 1907 23833 1916
rect 23885 1907 23904 1916
rect 23956 1907 23975 1916
rect 24027 1907 24046 1916
rect 24098 1910 24356 1916
rect 24098 1907 24104 1910
tri 24104 1907 24107 1910 nw
rect 22236 1865 22248 1875
rect 22282 1865 22288 1875
rect 22236 1863 22288 1865
rect 22236 1799 22248 1811
rect 22282 1799 22288 1811
tri 22430 1800 22433 1803 se
rect 22433 1800 22439 1803
rect 22354 1794 22439 1800
rect 22354 1760 22366 1794
rect 22400 1760 22438 1794
rect 22354 1754 22439 1760
tri 22430 1751 22433 1754 ne
rect 22433 1751 22439 1754
rect 22491 1751 22507 1803
rect 22559 1751 22575 1803
rect 22627 1751 22643 1803
rect 22695 1751 22711 1803
rect 22763 1751 22779 1803
rect 22831 1794 22847 1803
rect 22899 1794 22915 1803
rect 22967 1794 22982 1803
rect 23034 1794 23049 1803
rect 23101 1794 23116 1803
rect 23168 1794 23183 1803
rect 23235 1794 23250 1803
rect 23302 1800 23308 1803
tri 23308 1800 23311 1803 sw
rect 23302 1794 24356 1800
rect 22832 1760 22847 1794
rect 22904 1760 22915 1794
rect 22976 1760 22982 1794
rect 23048 1760 23049 1794
rect 23336 1760 23374 1794
rect 23408 1760 23446 1794
rect 23480 1760 23518 1794
rect 23552 1760 23590 1794
rect 23624 1760 23662 1794
rect 23696 1760 23734 1794
rect 23768 1760 23806 1794
rect 23840 1760 23878 1794
rect 23912 1760 23950 1794
rect 23984 1760 24022 1794
rect 24056 1760 24094 1794
rect 24128 1760 24166 1794
rect 24200 1760 24238 1794
rect 24272 1760 24310 1794
rect 24344 1760 24356 1794
rect 22831 1751 22847 1760
rect 22899 1751 22915 1760
rect 22967 1751 22982 1760
rect 23034 1751 23049 1760
rect 23101 1751 23116 1760
rect 23168 1751 23183 1760
rect 23235 1751 23250 1760
rect 23302 1754 24356 1760
rect 23302 1751 23308 1754
tri 23308 1751 23311 1754 nw
rect 22236 1735 22248 1747
rect 22282 1735 22288 1747
rect 22236 1672 22288 1683
rect 22236 1671 22248 1672
rect 22282 1671 22288 1672
tri 23398 1644 23401 1647 se
rect 23401 1644 23407 1647
rect 22236 1607 22288 1619
rect 22354 1638 23407 1644
rect 23459 1638 23478 1647
rect 23530 1638 23549 1647
rect 23601 1638 23620 1647
rect 23672 1638 23691 1647
rect 23743 1638 23762 1647
rect 23814 1638 23833 1647
rect 23885 1638 23904 1647
rect 23956 1638 23975 1647
rect 24027 1638 24046 1647
rect 24098 1644 24104 1647
tri 24104 1644 24107 1647 sw
rect 24098 1638 24356 1644
rect 22354 1604 22366 1638
rect 22400 1604 22438 1638
rect 22472 1604 22510 1638
rect 22544 1604 22582 1638
rect 22616 1604 22654 1638
rect 22688 1604 22726 1638
rect 22760 1604 22798 1638
rect 22832 1604 22870 1638
rect 22904 1604 22942 1638
rect 22976 1604 23014 1638
rect 23048 1604 23086 1638
rect 23120 1604 23158 1638
rect 23192 1604 23230 1638
rect 23264 1604 23302 1638
rect 23336 1604 23374 1638
rect 24128 1604 24166 1638
rect 24200 1604 24238 1638
rect 24272 1604 24310 1638
rect 24344 1604 24356 1638
rect 22354 1598 23407 1604
tri 23398 1595 23401 1598 ne
rect 23401 1595 23407 1598
rect 23459 1595 23478 1604
rect 23530 1595 23549 1604
rect 23601 1595 23620 1604
rect 23672 1595 23691 1604
rect 23743 1595 23762 1604
rect 23814 1595 23833 1604
rect 23885 1595 23904 1604
rect 23956 1595 23975 1604
rect 24027 1595 24046 1604
rect 24098 1598 24356 1604
rect 24098 1595 24104 1598
tri 24104 1595 24107 1598 nw
rect 22236 1543 22288 1555
rect 22236 1486 22248 1491
rect 22282 1486 22288 1491
tri 22430 1488 22433 1491 se
rect 22433 1488 22439 1491
rect 22236 1479 22288 1486
rect 22354 1482 22439 1488
rect 22354 1448 22366 1482
rect 22400 1448 22438 1482
rect 22354 1442 22439 1448
tri 22430 1439 22433 1442 ne
rect 22433 1439 22439 1442
rect 22491 1439 22507 1491
rect 22559 1439 22575 1491
rect 22627 1439 22643 1491
rect 22695 1439 22711 1491
rect 22763 1439 22779 1491
rect 22831 1482 22847 1491
rect 22899 1482 22915 1491
rect 22967 1482 22982 1491
rect 23034 1482 23049 1491
rect 23101 1482 23116 1491
rect 23168 1482 23183 1491
rect 23235 1482 23250 1491
rect 23302 1488 23308 1491
tri 23308 1488 23311 1491 sw
rect 23302 1482 24356 1488
rect 22832 1448 22847 1482
rect 22904 1448 22915 1482
rect 22976 1448 22982 1482
rect 23048 1448 23049 1482
rect 23336 1448 23374 1482
rect 23408 1448 23446 1482
rect 23480 1448 23518 1482
rect 23552 1448 23590 1482
rect 23624 1448 23662 1482
rect 23696 1448 23734 1482
rect 23768 1448 23806 1482
rect 23840 1448 23878 1482
rect 23912 1448 23950 1482
rect 23984 1448 24022 1482
rect 24056 1448 24094 1482
rect 24128 1448 24166 1482
rect 24200 1448 24238 1482
rect 24272 1448 24310 1482
rect 24344 1448 24356 1482
rect 22831 1439 22847 1448
rect 22899 1439 22915 1448
rect 22967 1439 22982 1448
rect 23034 1439 23049 1448
rect 23101 1439 23116 1448
rect 23168 1439 23183 1448
rect 23235 1439 23250 1448
rect 23302 1442 24356 1448
rect 23302 1439 23308 1442
tri 23308 1439 23311 1442 nw
rect 22236 1415 22248 1427
rect 22282 1415 22288 1427
rect 22236 1351 22248 1363
rect 22282 1351 22288 1363
tri 23398 1332 23401 1335 se
rect 23401 1332 23407 1335
rect 22236 1292 22288 1299
rect 22236 1287 22248 1292
rect 22282 1287 22288 1292
rect 7610 1266 7616 1269
rect 6371 1260 7616 1266
rect 7668 1260 7681 1269
rect 6371 1226 6383 1260
rect 6417 1226 6455 1260
rect 6489 1226 6527 1260
rect 6561 1226 6599 1260
rect 6633 1226 6671 1260
rect 6705 1226 6743 1260
rect 6777 1226 6815 1260
rect 6849 1226 6887 1260
rect 6921 1226 6959 1260
rect 6993 1226 7031 1260
rect 7065 1226 7103 1260
rect 7137 1226 7175 1260
rect 7209 1226 7247 1260
rect 7281 1226 7319 1260
rect 7353 1226 7391 1260
rect 7425 1226 7463 1260
rect 7497 1226 7535 1260
rect 7569 1226 7607 1260
rect 7668 1226 7679 1260
rect 6371 1220 7616 1226
rect 7610 1217 7616 1220
rect 7668 1217 7681 1226
rect 7733 1217 7746 1269
rect 7798 1217 7811 1269
rect 7863 1217 7876 1269
rect 7928 1260 7941 1269
rect 7993 1260 8006 1269
rect 8058 1260 8071 1269
rect 8123 1260 8136 1269
rect 8188 1260 8201 1269
rect 8253 1260 8266 1269
rect 8318 1260 8331 1269
rect 7929 1226 7941 1260
rect 8001 1226 8006 1260
rect 8253 1226 8255 1260
rect 8318 1226 8327 1260
rect 7928 1217 7941 1226
rect 7993 1217 8006 1226
rect 8058 1217 8071 1226
rect 8123 1217 8136 1226
rect 8188 1217 8201 1226
rect 8253 1217 8266 1226
rect 8318 1217 8331 1226
rect 8383 1217 8396 1269
rect 8448 1217 8461 1269
rect 8513 1217 8526 1269
rect 8578 1217 8591 1269
rect 8643 1260 8656 1269
rect 8708 1260 8721 1269
rect 8773 1260 8786 1269
rect 8838 1260 8851 1269
rect 8903 1260 8916 1269
rect 8968 1260 8981 1269
rect 8649 1226 8656 1260
rect 8968 1226 8975 1260
rect 8643 1217 8656 1226
rect 8708 1217 8721 1226
rect 8773 1217 8786 1226
rect 8838 1217 8851 1226
rect 8903 1217 8916 1226
rect 8968 1217 8981 1226
rect 9033 1217 9046 1269
rect 9098 1217 9111 1269
rect 9163 1217 9176 1269
rect 9228 1217 9241 1269
rect 9293 1260 9306 1269
rect 9358 1260 9371 1269
rect 9297 1226 9306 1260
rect 9369 1226 9371 1260
rect 9293 1217 9306 1226
rect 9358 1217 9371 1226
rect 9423 1217 9436 1269
rect 9488 1217 9501 1269
rect 9553 1260 9566 1269
rect 9618 1260 9631 1269
rect 9683 1260 9696 1269
rect 9748 1260 9761 1269
rect 9813 1260 9826 1269
rect 9748 1226 9749 1260
rect 9813 1226 9821 1260
rect 9553 1217 9566 1226
rect 9618 1217 9631 1226
rect 9683 1217 9696 1226
rect 9748 1217 9761 1226
rect 9813 1217 9826 1226
rect 9878 1217 9891 1269
rect 9943 1217 9956 1269
rect 10008 1217 10021 1269
rect 10073 1217 10086 1269
rect 10138 1260 10151 1269
rect 10203 1260 10216 1269
rect 10268 1260 10281 1269
rect 10333 1260 10346 1269
rect 10398 1260 10411 1269
rect 10463 1260 10476 1269
rect 10143 1226 10151 1260
rect 10215 1226 10216 1260
rect 10463 1226 10469 1260
rect 10138 1217 10151 1226
rect 10203 1217 10216 1226
rect 10268 1217 10281 1226
rect 10333 1217 10346 1226
rect 10398 1217 10411 1226
rect 10463 1217 10476 1226
rect 10528 1217 10541 1269
rect 10593 1217 10606 1269
rect 10658 1217 10671 1269
rect 10723 1217 10736 1269
rect 10788 1260 10800 1269
rect 10852 1260 10864 1269
rect 10916 1260 10928 1269
rect 10980 1260 10992 1269
rect 11044 1260 11056 1269
rect 11108 1260 11120 1269
rect 10791 1226 10800 1260
rect 10863 1226 10864 1260
rect 11044 1226 11045 1260
rect 11108 1226 11117 1260
rect 10788 1217 10800 1226
rect 10852 1217 10864 1226
rect 10916 1217 10928 1226
rect 10980 1217 10992 1226
rect 11044 1217 11056 1226
rect 11108 1217 11120 1226
rect 11172 1217 11184 1269
rect 11236 1217 11248 1269
rect 11300 1217 11312 1269
rect 11364 1260 11376 1269
rect 11428 1260 11440 1269
rect 11492 1260 11504 1269
rect 11556 1260 11568 1269
rect 11620 1260 11632 1269
rect 11684 1260 11696 1269
rect 11367 1226 11376 1260
rect 11439 1226 11440 1260
rect 11620 1226 11621 1260
rect 11684 1226 11693 1260
rect 11364 1217 11376 1226
rect 11428 1217 11440 1226
rect 11492 1217 11504 1226
rect 11556 1217 11568 1226
rect 11620 1217 11632 1226
rect 11684 1217 11696 1226
rect 11748 1217 11760 1269
rect 11812 1217 11824 1269
rect 11876 1266 11882 1269
rect 11876 1260 12531 1266
rect 11876 1226 11909 1260
rect 11943 1226 11981 1260
rect 12015 1226 12053 1260
rect 12087 1226 12125 1260
rect 12159 1226 12197 1260
rect 12231 1226 12269 1260
rect 12303 1226 12341 1260
rect 12375 1226 12413 1260
rect 12447 1226 12485 1260
rect 12519 1226 12531 1260
rect 11876 1220 12531 1226
rect 11876 1217 11882 1220
rect 12588 1218 12594 1270
rect 12646 1218 12659 1270
rect 12711 1260 12724 1270
rect 12776 1260 12789 1270
rect 12841 1260 12854 1270
rect 12906 1260 12919 1270
rect 12971 1260 12984 1270
rect 13036 1260 13049 1270
rect 12717 1226 12724 1260
rect 13036 1226 13043 1260
rect 12711 1218 12724 1226
rect 12776 1218 12789 1226
rect 12841 1218 12854 1226
rect 12906 1218 12919 1226
rect 12971 1218 12984 1226
rect 13036 1218 13049 1226
rect 13101 1218 13114 1270
rect 13166 1218 13179 1270
rect 13231 1218 13244 1270
rect 13296 1218 13309 1270
rect 13361 1260 13374 1270
rect 13426 1260 13439 1270
rect 13491 1260 13504 1270
rect 13556 1260 13569 1270
rect 13621 1260 13633 1270
rect 13685 1260 13697 1270
rect 13365 1226 13374 1260
rect 13437 1226 13439 1260
rect 13685 1226 13691 1260
rect 13361 1218 13374 1226
rect 13426 1218 13439 1226
rect 13491 1218 13504 1226
rect 13556 1218 13569 1226
rect 13621 1218 13633 1226
rect 13685 1218 13697 1226
rect 13749 1218 13761 1270
rect 13813 1218 13825 1270
rect 13877 1218 13889 1270
rect 13941 1218 13953 1270
rect 14005 1260 14017 1270
rect 14069 1260 14081 1270
rect 14133 1260 14145 1270
rect 14197 1260 14209 1270
rect 14261 1260 14273 1270
rect 14013 1226 14017 1260
rect 14261 1226 14267 1260
rect 14005 1218 14017 1226
rect 14069 1218 14081 1226
rect 14133 1218 14145 1226
rect 14197 1218 14209 1226
rect 14261 1218 14273 1226
rect 14325 1218 14337 1270
rect 14389 1218 14401 1270
rect 14453 1218 14465 1270
rect 14517 1218 14529 1270
rect 14581 1260 14593 1270
rect 14645 1260 14657 1270
rect 14709 1260 14721 1270
rect 14773 1260 14785 1270
rect 14837 1260 14849 1270
rect 14589 1226 14593 1260
rect 14837 1226 14843 1260
rect 14581 1218 14593 1226
rect 14645 1218 14657 1226
rect 14709 1218 14721 1226
rect 14773 1218 14785 1226
rect 14837 1218 14849 1226
rect 14901 1218 14913 1270
rect 14965 1218 14977 1270
rect 15029 1218 15041 1270
rect 15093 1218 15105 1270
rect 15157 1260 15169 1270
rect 15221 1260 15233 1270
rect 15285 1260 15297 1270
rect 15349 1260 15361 1270
rect 15413 1260 15425 1270
rect 15165 1226 15169 1260
rect 15413 1226 15419 1260
rect 15157 1218 15169 1226
rect 15221 1218 15233 1226
rect 15285 1218 15297 1226
rect 15349 1218 15361 1226
rect 15413 1218 15425 1226
rect 15477 1218 15489 1270
rect 15541 1218 15553 1270
rect 15605 1218 15617 1270
rect 15669 1218 15681 1270
rect 15733 1218 15745 1270
rect 15797 1218 15809 1270
rect 15861 1260 15873 1270
rect 15925 1260 15937 1270
rect 15989 1260 16001 1270
rect 16053 1260 16065 1270
rect 16117 1260 16129 1270
rect 15867 1226 15873 1260
rect 16117 1226 16121 1260
rect 15861 1218 15873 1226
rect 15925 1218 15937 1226
rect 15989 1218 16001 1226
rect 16053 1218 16065 1226
rect 16117 1218 16129 1226
rect 16181 1218 16193 1270
rect 16245 1218 16257 1270
rect 16309 1218 16321 1270
rect 16373 1218 16385 1270
rect 16437 1260 16449 1270
rect 16501 1260 16513 1270
rect 16565 1260 16577 1270
rect 16629 1260 16641 1270
rect 16693 1260 16705 1270
rect 16443 1226 16449 1260
rect 16693 1226 16697 1260
rect 16437 1218 16449 1226
rect 16501 1218 16513 1226
rect 16565 1218 16577 1226
rect 16629 1218 16641 1226
rect 16693 1218 16705 1226
rect 16757 1218 16769 1270
rect 16821 1218 16833 1270
rect 16885 1218 16897 1270
rect 16949 1218 16961 1270
rect 17013 1260 17025 1270
rect 17077 1260 17089 1270
rect 17141 1260 17153 1270
rect 17205 1260 17217 1270
rect 17269 1260 17281 1270
rect 17019 1226 17025 1260
rect 17269 1226 17273 1260
rect 17013 1218 17025 1226
rect 17077 1218 17089 1226
rect 17141 1218 17153 1226
rect 17205 1218 17217 1226
rect 17269 1218 17281 1226
rect 17333 1218 17345 1270
rect 17397 1218 17409 1270
rect 17461 1218 17473 1270
rect 17525 1218 17537 1270
rect 17589 1260 17601 1270
rect 17653 1260 17665 1270
rect 17717 1260 17729 1270
rect 17781 1260 17793 1270
rect 17845 1260 17857 1270
rect 17595 1226 17601 1260
rect 17845 1226 17849 1260
rect 17589 1218 17601 1226
rect 17653 1218 17665 1226
rect 17717 1218 17729 1226
rect 17781 1218 17793 1226
rect 17845 1218 17857 1226
rect 17909 1218 17921 1270
rect 17973 1218 17985 1270
rect 18037 1218 18049 1270
rect 18101 1218 18113 1270
rect 18165 1260 18177 1270
rect 18229 1260 18241 1270
rect 18293 1260 18305 1270
rect 18357 1260 18369 1270
rect 18421 1260 18433 1270
rect 18171 1226 18177 1260
rect 18421 1226 18425 1260
rect 18165 1218 18177 1226
rect 18229 1218 18241 1226
rect 18293 1218 18305 1226
rect 18357 1218 18369 1226
rect 18421 1218 18433 1226
rect 18485 1218 18497 1270
rect 18549 1218 18561 1270
rect 18613 1218 18625 1270
rect 18677 1218 18689 1270
rect 18741 1260 18753 1270
rect 18805 1260 18817 1270
rect 18747 1226 18753 1260
rect 18741 1218 18753 1226
rect 18805 1218 18817 1226
rect 18869 1218 18881 1270
rect 18933 1218 18945 1270
rect 18997 1260 19009 1270
rect 19061 1260 19073 1270
rect 19125 1260 19137 1270
rect 19189 1260 19201 1270
rect 19125 1226 19127 1260
rect 19189 1226 19199 1260
rect 18997 1218 19009 1226
rect 19061 1218 19073 1226
rect 19125 1218 19137 1226
rect 19189 1218 19201 1226
rect 19253 1218 19265 1270
rect 19317 1218 19329 1270
rect 19381 1218 19393 1270
rect 19445 1260 19457 1270
rect 19509 1260 19521 1270
rect 19573 1260 19585 1270
rect 19637 1260 19649 1270
rect 19701 1260 19713 1270
rect 19765 1260 19777 1270
rect 19449 1226 19457 1260
rect 19701 1226 19703 1260
rect 19765 1226 19775 1260
rect 19445 1218 19457 1226
rect 19509 1218 19521 1226
rect 19573 1218 19585 1226
rect 19637 1218 19649 1226
rect 19701 1218 19713 1226
rect 19765 1218 19777 1226
rect 19829 1218 19841 1270
rect 19893 1218 19905 1270
rect 19957 1218 19969 1270
rect 20021 1260 20033 1270
rect 20085 1260 20097 1270
rect 20149 1260 20161 1270
rect 20213 1260 20225 1270
rect 20277 1260 20289 1270
rect 20341 1260 20353 1270
rect 20025 1226 20033 1260
rect 20277 1226 20279 1260
rect 20341 1226 20351 1260
rect 20021 1218 20033 1226
rect 20085 1218 20097 1226
rect 20149 1218 20161 1226
rect 20213 1218 20225 1226
rect 20277 1218 20289 1226
rect 20341 1218 20353 1226
rect 20405 1218 20417 1270
rect 20469 1218 20481 1270
rect 20533 1218 20545 1270
rect 20597 1260 20609 1270
rect 20661 1260 20673 1270
rect 20725 1260 20737 1270
rect 20789 1260 20801 1270
rect 20853 1260 20865 1270
rect 20917 1260 20929 1270
rect 20601 1226 20609 1260
rect 20853 1226 20855 1260
rect 20917 1226 20927 1260
rect 20597 1218 20609 1226
rect 20661 1218 20673 1226
rect 20725 1218 20737 1226
rect 20789 1218 20801 1226
rect 20853 1218 20865 1226
rect 20917 1218 20929 1226
rect 20981 1218 20993 1270
rect 21045 1218 21057 1270
rect 21109 1218 21121 1270
rect 21173 1260 21185 1270
rect 21237 1260 21249 1270
rect 21301 1260 21313 1270
rect 21365 1260 21377 1270
rect 21429 1260 21441 1270
rect 21493 1260 21505 1270
rect 21177 1226 21185 1260
rect 21429 1226 21431 1260
rect 21493 1226 21503 1260
rect 21173 1218 21185 1226
rect 21237 1218 21249 1226
rect 21301 1218 21313 1226
rect 21365 1218 21377 1226
rect 21429 1218 21441 1226
rect 21493 1218 21505 1226
rect 21557 1218 21569 1270
rect 21621 1218 21633 1270
rect 21685 1218 21697 1270
rect 21749 1260 21761 1270
rect 21813 1260 21825 1270
rect 21877 1260 21889 1270
rect 21941 1266 21947 1270
rect 21941 1260 21981 1266
rect 21753 1226 21761 1260
rect 21969 1226 21981 1260
rect 21749 1218 21761 1226
rect 21813 1218 21825 1226
rect 21877 1218 21889 1226
rect 21941 1220 21981 1226
rect 22354 1326 23407 1332
rect 23459 1326 23478 1335
rect 23530 1326 23549 1335
rect 23601 1326 23620 1335
rect 23672 1326 23691 1335
rect 23743 1326 23762 1335
rect 23814 1326 23833 1335
rect 23885 1326 23904 1335
rect 23956 1326 23975 1335
rect 24027 1326 24046 1335
rect 24098 1332 24104 1335
tri 24104 1332 24107 1335 sw
rect 24098 1326 24356 1332
rect 22354 1292 22366 1326
rect 22400 1292 22438 1326
rect 22472 1292 22510 1326
rect 22544 1292 22582 1326
rect 22616 1292 22654 1326
rect 22688 1292 22726 1326
rect 22760 1292 22798 1326
rect 22832 1292 22870 1326
rect 22904 1292 22942 1326
rect 22976 1292 23014 1326
rect 23048 1292 23086 1326
rect 23120 1292 23158 1326
rect 23192 1292 23230 1326
rect 23264 1292 23302 1326
rect 23336 1292 23374 1326
rect 24128 1292 24166 1326
rect 24200 1292 24238 1326
rect 24272 1292 24310 1326
rect 24344 1292 24356 1326
rect 22354 1286 23407 1292
tri 23398 1283 23401 1286 ne
rect 23401 1283 23407 1286
rect 23459 1283 23478 1292
rect 23530 1283 23549 1292
rect 23601 1283 23620 1292
rect 23672 1283 23691 1292
rect 23743 1283 23762 1292
rect 23814 1283 23833 1292
rect 23885 1283 23904 1292
rect 23956 1283 23975 1292
rect 24027 1283 24046 1292
rect 24098 1286 24356 1292
rect 24098 1283 24104 1286
tri 24104 1283 24107 1286 nw
rect 22236 1223 22288 1235
rect 21941 1218 21947 1220
rect 6267 1183 22236 1189
rect 6267 1177 9388 1183
rect 6267 1143 6273 1177
rect 6307 1149 9388 1177
rect 9422 1149 9460 1183
rect 9494 1149 12538 1183
rect 12572 1149 12610 1183
rect 12644 1149 15688 1183
rect 15722 1149 15760 1183
rect 15794 1149 18838 1183
rect 18872 1149 18910 1183
rect 18944 1149 21988 1183
rect 22022 1149 22060 1183
rect 22094 1171 22236 1183
tri 22430 1176 22433 1179 se
rect 22433 1176 22439 1179
rect 22094 1159 22288 1171
rect 22094 1149 22236 1159
rect 6307 1143 22236 1149
rect 6267 1140 6337 1143
tri 6337 1140 6340 1143 nw
rect 6267 1102 6313 1140
tri 6313 1116 6337 1140 nw
rect 7610 1110 7616 1113
rect 6267 1068 6273 1102
rect 6307 1068 6313 1102
rect 6267 1033 6313 1068
rect 6371 1104 7616 1110
rect 7668 1104 7681 1113
rect 6371 1070 6383 1104
rect 6417 1070 6455 1104
rect 6489 1070 6527 1104
rect 6561 1070 6599 1104
rect 6633 1070 6671 1104
rect 6705 1070 6743 1104
rect 6777 1070 6815 1104
rect 6849 1070 6887 1104
rect 6921 1070 6959 1104
rect 6993 1070 7031 1104
rect 7065 1070 7103 1104
rect 7137 1070 7175 1104
rect 7209 1070 7247 1104
rect 7281 1070 7319 1104
rect 7353 1070 7391 1104
rect 7425 1070 7463 1104
rect 7497 1070 7535 1104
rect 7569 1070 7607 1104
rect 7668 1070 7679 1104
rect 6371 1064 7616 1070
rect 7610 1061 7616 1064
rect 7668 1061 7681 1070
rect 7733 1061 7746 1113
rect 7798 1061 7811 1113
rect 7863 1061 7876 1113
rect 7928 1104 7941 1113
rect 7993 1104 8006 1113
rect 8058 1104 8071 1113
rect 8123 1104 8136 1113
rect 8188 1104 8201 1113
rect 8253 1104 8266 1113
rect 8318 1104 8331 1113
rect 7929 1070 7941 1104
rect 8001 1070 8006 1104
rect 8253 1070 8255 1104
rect 8318 1070 8327 1104
rect 7928 1061 7941 1070
rect 7993 1061 8006 1070
rect 8058 1061 8071 1070
rect 8123 1061 8136 1070
rect 8188 1061 8201 1070
rect 8253 1061 8266 1070
rect 8318 1061 8331 1070
rect 8383 1061 8396 1113
rect 8448 1061 8461 1113
rect 8513 1061 8526 1113
rect 8578 1061 8591 1113
rect 8643 1104 8656 1113
rect 8708 1104 8721 1113
rect 8773 1104 8786 1113
rect 8838 1104 8851 1113
rect 8903 1104 8916 1113
rect 8968 1104 8981 1113
rect 8649 1070 8656 1104
rect 8968 1070 8975 1104
rect 8643 1061 8656 1070
rect 8708 1061 8721 1070
rect 8773 1061 8786 1070
rect 8838 1061 8851 1070
rect 8903 1061 8916 1070
rect 8968 1061 8981 1070
rect 9033 1061 9046 1113
rect 9098 1061 9111 1113
rect 9163 1061 9176 1113
rect 9228 1061 9241 1113
rect 9293 1104 9306 1113
rect 9358 1104 9371 1113
rect 9297 1070 9306 1104
rect 9369 1070 9371 1104
rect 9293 1061 9306 1070
rect 9358 1061 9371 1070
rect 9423 1061 9436 1113
rect 9488 1061 9501 1113
rect 9553 1104 9566 1113
rect 9618 1104 9631 1113
rect 9683 1104 9696 1113
rect 9748 1104 9761 1113
rect 9813 1104 9826 1113
rect 9748 1070 9749 1104
rect 9813 1070 9821 1104
rect 9553 1061 9566 1070
rect 9618 1061 9631 1070
rect 9683 1061 9696 1070
rect 9748 1061 9761 1070
rect 9813 1061 9826 1070
rect 9878 1061 9891 1113
rect 9943 1061 9956 1113
rect 10008 1061 10021 1113
rect 10073 1061 10086 1113
rect 10138 1104 10151 1113
rect 10203 1104 10216 1113
rect 10268 1104 10281 1113
rect 10333 1104 10346 1113
rect 10398 1104 10411 1113
rect 10463 1104 10476 1113
rect 10143 1070 10151 1104
rect 10215 1070 10216 1104
rect 10463 1070 10469 1104
rect 10138 1061 10151 1070
rect 10203 1061 10216 1070
rect 10268 1061 10281 1070
rect 10333 1061 10346 1070
rect 10398 1061 10411 1070
rect 10463 1061 10476 1070
rect 10528 1061 10541 1113
rect 10593 1061 10606 1113
rect 10658 1061 10671 1113
rect 10723 1061 10736 1113
rect 10788 1104 10800 1113
rect 10852 1104 10864 1113
rect 10916 1104 10928 1113
rect 10980 1104 10992 1113
rect 11044 1104 11056 1113
rect 11108 1104 11120 1113
rect 10791 1070 10800 1104
rect 10863 1070 10864 1104
rect 11044 1070 11045 1104
rect 11108 1070 11117 1104
rect 10788 1061 10800 1070
rect 10852 1061 10864 1070
rect 10916 1061 10928 1070
rect 10980 1061 10992 1070
rect 11044 1061 11056 1070
rect 11108 1061 11120 1070
rect 11172 1061 11184 1113
rect 11236 1061 11248 1113
rect 11300 1061 11312 1113
rect 11364 1104 11376 1113
rect 11428 1104 11440 1113
rect 11492 1104 11504 1113
rect 11556 1104 11568 1113
rect 11620 1104 11632 1113
rect 11684 1104 11696 1113
rect 11367 1070 11376 1104
rect 11439 1070 11440 1104
rect 11620 1070 11621 1104
rect 11684 1070 11693 1104
rect 11364 1061 11376 1070
rect 11428 1061 11440 1070
rect 11492 1061 11504 1070
rect 11556 1061 11568 1070
rect 11620 1061 11632 1070
rect 11684 1061 11696 1070
rect 11748 1061 11760 1113
rect 11812 1061 11824 1113
rect 11876 1110 11882 1113
rect 12016 1110 12022 1113
rect 11876 1104 12022 1110
rect 12074 1104 12087 1113
rect 12139 1104 12152 1113
rect 12204 1104 12217 1113
rect 12269 1104 12282 1113
rect 12334 1104 12347 1113
rect 11876 1070 11909 1104
rect 11943 1070 11981 1104
rect 12015 1070 12022 1104
rect 12334 1070 12341 1104
rect 11876 1064 12022 1070
rect 11876 1061 11882 1064
rect 12016 1061 12022 1064
rect 12074 1061 12087 1070
rect 12139 1061 12152 1070
rect 12204 1061 12217 1070
rect 12269 1061 12282 1070
rect 12334 1061 12347 1070
rect 12399 1061 12412 1113
rect 12464 1061 12477 1113
rect 12529 1061 12542 1113
rect 12594 1061 12607 1113
rect 12659 1061 12672 1113
rect 12724 1061 12737 1113
rect 12789 1061 12801 1113
rect 12853 1104 12865 1113
rect 12917 1104 12929 1113
rect 12981 1104 12993 1113
rect 13045 1104 13057 1113
rect 13109 1104 13121 1113
rect 12861 1070 12865 1104
rect 13109 1070 13115 1104
rect 12853 1061 12865 1070
rect 12917 1061 12929 1070
rect 12981 1061 12993 1070
rect 13045 1061 13057 1070
rect 13109 1061 13121 1070
rect 13173 1061 13185 1113
rect 13237 1061 13249 1113
rect 13301 1061 13313 1113
rect 13365 1061 13377 1113
rect 13429 1104 13441 1113
rect 13493 1104 13505 1113
rect 13557 1104 13569 1113
rect 13621 1104 13633 1113
rect 13685 1104 13697 1113
rect 13437 1070 13441 1104
rect 13685 1070 13691 1104
rect 13429 1061 13441 1070
rect 13493 1061 13505 1070
rect 13557 1061 13569 1070
rect 13621 1061 13633 1070
rect 13685 1061 13697 1070
rect 13749 1061 13761 1113
rect 13813 1061 13825 1113
rect 13877 1061 13889 1113
rect 13941 1061 13953 1113
rect 14005 1104 14017 1113
rect 14069 1104 14081 1113
rect 14133 1104 14145 1113
rect 14197 1104 14209 1113
rect 14261 1104 14273 1113
rect 14013 1070 14017 1104
rect 14261 1070 14267 1104
rect 14005 1061 14017 1070
rect 14069 1061 14081 1070
rect 14133 1061 14145 1070
rect 14197 1061 14209 1070
rect 14261 1061 14273 1070
rect 14325 1061 14337 1113
rect 14389 1061 14401 1113
rect 14453 1061 14465 1113
rect 14517 1061 14529 1113
rect 14581 1104 14593 1113
rect 14645 1104 14657 1113
rect 14709 1104 14721 1113
rect 14773 1104 14785 1113
rect 14837 1104 14849 1113
rect 14589 1070 14593 1104
rect 14837 1070 14843 1104
rect 14581 1061 14593 1070
rect 14645 1061 14657 1070
rect 14709 1061 14721 1070
rect 14773 1061 14785 1070
rect 14837 1061 14849 1070
rect 14901 1061 14913 1113
rect 14965 1061 14977 1113
rect 15029 1061 15041 1113
rect 15093 1061 15105 1113
rect 15157 1104 15169 1113
rect 15221 1104 15233 1113
rect 15285 1104 15297 1113
rect 15349 1104 15361 1113
rect 15413 1104 15425 1113
rect 15165 1070 15169 1104
rect 15413 1070 15419 1104
rect 15157 1061 15169 1070
rect 15221 1061 15233 1070
rect 15285 1061 15297 1070
rect 15349 1061 15361 1070
rect 15413 1061 15425 1070
rect 15477 1061 15489 1113
rect 15541 1061 15553 1113
rect 15605 1061 15617 1113
rect 15669 1061 15681 1113
rect 15733 1061 15745 1113
rect 15797 1061 15809 1113
rect 15861 1104 15873 1113
rect 15925 1104 15937 1113
rect 15989 1104 16001 1113
rect 16053 1104 16065 1113
rect 16117 1104 16129 1113
rect 15867 1070 15873 1104
rect 16117 1070 16121 1104
rect 15861 1061 15873 1070
rect 15925 1061 15937 1070
rect 15989 1061 16001 1070
rect 16053 1061 16065 1070
rect 16117 1061 16129 1070
rect 16181 1061 16193 1113
rect 16245 1061 16257 1113
rect 16309 1061 16321 1113
rect 16373 1061 16385 1113
rect 16437 1104 16449 1113
rect 16501 1104 16513 1113
rect 16565 1104 16577 1113
rect 16629 1104 16641 1113
rect 16693 1104 16705 1113
rect 16443 1070 16449 1104
rect 16693 1070 16697 1104
rect 16437 1061 16449 1070
rect 16501 1061 16513 1070
rect 16565 1061 16577 1070
rect 16629 1061 16641 1070
rect 16693 1061 16705 1070
rect 16757 1061 16769 1113
rect 16821 1061 16833 1113
rect 16885 1061 16897 1113
rect 16949 1061 16961 1113
rect 17013 1104 17025 1113
rect 17077 1104 17089 1113
rect 17141 1104 17153 1113
rect 17205 1104 17217 1113
rect 17269 1104 17281 1113
rect 17019 1070 17025 1104
rect 17269 1070 17273 1104
rect 17013 1061 17025 1070
rect 17077 1061 17089 1070
rect 17141 1061 17153 1070
rect 17205 1061 17217 1070
rect 17269 1061 17281 1070
rect 17333 1061 17345 1113
rect 17397 1061 17409 1113
rect 17461 1061 17473 1113
rect 17525 1061 17537 1113
rect 17589 1104 17601 1113
rect 17653 1104 17665 1113
rect 17717 1104 17729 1113
rect 17781 1104 17793 1113
rect 17845 1104 17857 1113
rect 17595 1070 17601 1104
rect 17845 1070 17849 1104
rect 17589 1061 17601 1070
rect 17653 1061 17665 1070
rect 17717 1061 17729 1070
rect 17781 1061 17793 1070
rect 17845 1061 17857 1070
rect 17909 1061 17921 1113
rect 17973 1061 17985 1113
rect 18037 1061 18049 1113
rect 18101 1061 18113 1113
rect 18165 1104 18177 1113
rect 18229 1104 18241 1113
rect 18293 1104 18305 1113
rect 18357 1104 18369 1113
rect 18421 1104 18433 1113
rect 18171 1070 18177 1104
rect 18421 1070 18425 1104
rect 18165 1061 18177 1070
rect 18229 1061 18241 1070
rect 18293 1061 18305 1070
rect 18357 1061 18369 1070
rect 18421 1061 18433 1070
rect 18485 1061 18497 1113
rect 18549 1061 18561 1113
rect 18613 1061 18625 1113
rect 18677 1061 18689 1113
rect 18741 1104 18753 1113
rect 18805 1104 18817 1113
rect 18747 1070 18753 1104
rect 18741 1061 18753 1070
rect 18805 1061 18817 1070
rect 18869 1061 18881 1113
rect 18933 1061 18945 1113
rect 18997 1104 19009 1113
rect 19061 1104 19073 1113
rect 19125 1104 19137 1113
rect 19189 1104 19201 1113
rect 19125 1070 19127 1104
rect 19189 1070 19199 1104
rect 18997 1061 19009 1070
rect 19061 1061 19073 1070
rect 19125 1061 19137 1070
rect 19189 1061 19201 1070
rect 19253 1061 19265 1113
rect 19317 1061 19329 1113
rect 19381 1061 19393 1113
rect 19445 1104 19457 1113
rect 19509 1104 19521 1113
rect 19573 1104 19585 1113
rect 19637 1104 19649 1113
rect 19701 1104 19713 1113
rect 19765 1104 19777 1113
rect 19449 1070 19457 1104
rect 19701 1070 19703 1104
rect 19765 1070 19775 1104
rect 19445 1061 19457 1070
rect 19509 1061 19521 1070
rect 19573 1061 19585 1070
rect 19637 1061 19649 1070
rect 19701 1061 19713 1070
rect 19765 1061 19777 1070
rect 19829 1061 19841 1113
rect 19893 1061 19905 1113
rect 19957 1061 19969 1113
rect 20021 1104 20033 1113
rect 20085 1104 20097 1113
rect 20149 1104 20161 1113
rect 20213 1104 20225 1113
rect 20277 1104 20289 1113
rect 20341 1104 20353 1113
rect 20025 1070 20033 1104
rect 20277 1070 20279 1104
rect 20341 1070 20351 1104
rect 20021 1061 20033 1070
rect 20085 1061 20097 1070
rect 20149 1061 20161 1070
rect 20213 1061 20225 1070
rect 20277 1061 20289 1070
rect 20341 1061 20353 1070
rect 20405 1061 20417 1113
rect 20469 1061 20481 1113
rect 20533 1061 20545 1113
rect 20597 1104 20609 1113
rect 20661 1104 20673 1113
rect 20725 1104 20737 1113
rect 20789 1104 20801 1113
rect 20853 1104 20865 1113
rect 20917 1104 20929 1113
rect 20601 1070 20609 1104
rect 20853 1070 20855 1104
rect 20917 1070 20927 1104
rect 20597 1061 20609 1070
rect 20661 1061 20673 1070
rect 20725 1061 20737 1070
rect 20789 1061 20801 1070
rect 20853 1061 20865 1070
rect 20917 1061 20929 1070
rect 20981 1061 20993 1113
rect 21045 1061 21057 1113
rect 21109 1061 21121 1113
rect 21173 1104 21185 1113
rect 21237 1104 21249 1113
rect 21301 1104 21313 1113
rect 21365 1104 21377 1113
rect 21429 1104 21441 1113
rect 21493 1104 21505 1113
rect 21177 1070 21185 1104
rect 21429 1070 21431 1104
rect 21493 1070 21503 1104
rect 21173 1061 21185 1070
rect 21237 1061 21249 1070
rect 21301 1061 21313 1070
rect 21365 1061 21377 1070
rect 21429 1061 21441 1070
rect 21493 1061 21505 1070
rect 21557 1061 21569 1113
rect 21621 1061 21633 1113
rect 21685 1061 21697 1113
rect 21749 1104 21761 1113
rect 21813 1104 21825 1113
rect 21877 1104 21889 1113
rect 21941 1104 21981 1113
rect 21753 1070 21761 1104
rect 21969 1070 21981 1104
rect 21749 1061 21761 1070
rect 21813 1061 21825 1070
rect 21877 1061 21889 1070
rect 21941 1061 21981 1070
rect 22354 1170 22439 1176
rect 22354 1136 22366 1170
rect 22400 1136 22438 1170
rect 22354 1130 22439 1136
tri 22430 1127 22433 1130 ne
rect 22433 1127 22439 1130
rect 22491 1127 22507 1179
rect 22559 1127 22575 1179
rect 22627 1127 22643 1179
rect 22695 1127 22711 1179
rect 22763 1127 22779 1179
rect 22831 1170 22847 1179
rect 22899 1170 22915 1179
rect 22967 1170 22982 1179
rect 23034 1170 23049 1179
rect 23101 1170 23116 1179
rect 23168 1170 23183 1179
rect 23235 1170 23250 1179
rect 23302 1176 23308 1179
tri 23308 1176 23311 1179 sw
rect 23302 1170 24356 1176
rect 22832 1136 22847 1170
rect 22904 1136 22915 1170
rect 22976 1136 22982 1170
rect 23048 1136 23049 1170
rect 23336 1136 23374 1170
rect 23408 1136 23446 1170
rect 23480 1136 23518 1170
rect 23552 1136 23590 1170
rect 23624 1136 23662 1170
rect 23696 1136 23734 1170
rect 23768 1136 23806 1170
rect 23840 1136 23878 1170
rect 23912 1136 23950 1170
rect 23984 1136 24022 1170
rect 24056 1136 24094 1170
rect 24128 1136 24166 1170
rect 24200 1136 24238 1170
rect 24272 1136 24310 1170
rect 24344 1136 24356 1170
rect 22831 1127 22847 1136
rect 22899 1127 22915 1136
rect 22967 1127 22982 1136
rect 23034 1127 23049 1136
rect 23101 1127 23116 1136
rect 23168 1127 23183 1136
rect 23235 1127 23250 1136
rect 23302 1130 24356 1136
rect 23302 1127 23308 1130
tri 23308 1127 23311 1130 nw
rect 22236 1106 22248 1107
rect 22282 1106 22288 1107
rect 22236 1095 22288 1106
tri 6313 1033 6340 1060 sw
rect 22236 1033 22248 1043
rect 6267 1031 22248 1033
rect 22282 1031 22288 1043
rect 6267 1027 22236 1031
rect 6267 993 6273 1027
rect 6307 993 9388 1027
rect 9422 993 9460 1027
rect 9494 993 12538 1027
rect 12572 993 12610 1027
rect 12644 993 15688 1027
rect 15722 993 15760 1027
rect 15794 993 18838 1027
rect 18872 993 18910 1027
rect 18944 993 21988 1027
rect 22022 993 22060 1027
rect 22094 993 22236 1027
rect 6267 987 22236 993
tri 23399 1020 23401 1022 se
rect 23401 1020 23407 1022
rect 6267 952 6313 987
tri 6313 960 6340 987 nw
rect 22236 967 22248 979
rect 22282 967 22288 979
rect 22354 1014 23407 1020
rect 23459 1014 23478 1022
rect 23530 1014 23549 1022
rect 23601 1014 23620 1022
rect 23672 1014 23691 1022
rect 23743 1014 23762 1022
rect 23814 1014 23833 1022
rect 23885 1014 23904 1022
rect 23956 1014 23975 1022
rect 24027 1014 24046 1022
rect 24098 1020 24104 1022
tri 24104 1020 24106 1022 sw
rect 24098 1014 24356 1020
rect 22354 980 22366 1014
rect 22400 980 22438 1014
rect 22472 980 22510 1014
rect 22544 980 22582 1014
rect 22616 980 22654 1014
rect 22688 980 22726 1014
rect 22760 980 22798 1014
rect 22832 980 22870 1014
rect 22904 980 22942 1014
rect 22976 980 23014 1014
rect 23048 980 23086 1014
rect 23120 980 23158 1014
rect 23192 980 23230 1014
rect 23264 980 23302 1014
rect 23336 980 23374 1014
rect 24128 980 24166 1014
rect 24200 980 24238 1014
rect 24272 980 24310 1014
rect 24344 980 24356 1014
rect 22354 974 23407 980
tri 23397 970 23401 974 ne
rect 23401 970 23407 974
rect 23459 970 23478 980
rect 23530 970 23549 980
rect 23601 970 23620 980
rect 23672 970 23691 980
rect 23743 970 23762 980
rect 23814 970 23833 980
rect 23885 970 23904 980
rect 23956 970 23975 980
rect 24027 970 24046 980
rect 24098 974 24356 980
rect 24098 970 24104 974
tri 24104 970 24108 974 nw
rect 7610 954 7616 957
rect 6267 918 6273 952
rect 6307 918 6313 952
rect 6267 878 6313 918
rect 6371 948 7616 954
rect 7668 948 7681 957
rect 6371 914 6383 948
rect 6417 914 6455 948
rect 6489 914 6527 948
rect 6561 914 6599 948
rect 6633 914 6671 948
rect 6705 914 6743 948
rect 6777 914 6815 948
rect 6849 914 6887 948
rect 6921 914 6959 948
rect 6993 914 7031 948
rect 7065 914 7103 948
rect 7137 914 7175 948
rect 7209 914 7247 948
rect 7281 914 7319 948
rect 7353 914 7391 948
rect 7425 914 7463 948
rect 7497 914 7535 948
rect 7569 914 7607 948
rect 7668 914 7679 948
rect 6371 908 7616 914
rect 7610 905 7616 908
rect 7668 905 7681 914
rect 7733 905 7746 957
rect 7798 905 7811 957
rect 7863 905 7876 957
rect 7928 948 7941 957
rect 7993 948 8006 957
rect 8058 948 8071 957
rect 8123 948 8136 957
rect 8188 948 8201 957
rect 8253 948 8266 957
rect 8318 948 8331 957
rect 7929 914 7941 948
rect 8001 914 8006 948
rect 8253 914 8255 948
rect 8318 914 8327 948
rect 7928 905 7941 914
rect 7993 905 8006 914
rect 8058 905 8071 914
rect 8123 905 8136 914
rect 8188 905 8201 914
rect 8253 905 8266 914
rect 8318 905 8331 914
rect 8383 905 8396 957
rect 8448 905 8461 957
rect 8513 905 8526 957
rect 8578 905 8591 957
rect 8643 948 8656 957
rect 8708 948 8721 957
rect 8773 948 8786 957
rect 8838 948 8851 957
rect 8903 948 8916 957
rect 8968 948 8981 957
rect 8649 914 8656 948
rect 8968 914 8975 948
rect 8643 905 8656 914
rect 8708 905 8721 914
rect 8773 905 8786 914
rect 8838 905 8851 914
rect 8903 905 8916 914
rect 8968 905 8981 914
rect 9033 905 9046 957
rect 9098 905 9111 957
rect 9163 905 9176 957
rect 9228 905 9241 957
rect 9293 948 9306 957
rect 9358 948 9371 957
rect 9297 914 9306 948
rect 9369 914 9371 948
rect 9293 905 9306 914
rect 9358 905 9371 914
rect 9423 905 9436 957
rect 9488 905 9501 957
rect 9553 948 9566 957
rect 9618 948 9631 957
rect 9683 948 9696 957
rect 9748 948 9761 957
rect 9813 948 9826 957
rect 9748 914 9749 948
rect 9813 914 9821 948
rect 9553 905 9566 914
rect 9618 905 9631 914
rect 9683 905 9696 914
rect 9748 905 9761 914
rect 9813 905 9826 914
rect 9878 905 9891 957
rect 9943 905 9956 957
rect 10008 905 10021 957
rect 10073 905 10086 957
rect 10138 948 10151 957
rect 10203 948 10216 957
rect 10268 948 10281 957
rect 10333 948 10346 957
rect 10398 948 10411 957
rect 10463 948 10476 957
rect 10143 914 10151 948
rect 10215 914 10216 948
rect 10463 914 10469 948
rect 10138 905 10151 914
rect 10203 905 10216 914
rect 10268 905 10281 914
rect 10333 905 10346 914
rect 10398 905 10411 914
rect 10463 905 10476 914
rect 10528 905 10541 957
rect 10593 905 10606 957
rect 10658 905 10671 957
rect 10723 905 10736 957
rect 10788 948 10800 957
rect 10852 948 10864 957
rect 10916 948 10928 957
rect 10980 948 10992 957
rect 11044 948 11056 957
rect 11108 948 11120 957
rect 10791 914 10800 948
rect 10863 914 10864 948
rect 11044 914 11045 948
rect 11108 914 11117 948
rect 10788 905 10800 914
rect 10852 905 10864 914
rect 10916 905 10928 914
rect 10980 905 10992 914
rect 11044 905 11056 914
rect 11108 905 11120 914
rect 11172 905 11184 957
rect 11236 905 11248 957
rect 11300 905 11312 957
rect 11364 948 11376 957
rect 11428 948 11440 957
rect 11492 948 11504 957
rect 11556 948 11568 957
rect 11620 948 11632 957
rect 11684 948 11696 957
rect 11367 914 11376 948
rect 11439 914 11440 948
rect 11620 914 11621 948
rect 11684 914 11693 948
rect 11364 905 11376 914
rect 11428 905 11440 914
rect 11492 905 11504 914
rect 11556 905 11568 914
rect 11620 905 11632 914
rect 11684 905 11696 914
rect 11748 905 11760 957
rect 11812 905 11824 957
rect 11876 954 11882 957
rect 12016 954 12022 957
rect 11876 948 12022 954
rect 12074 948 12087 957
rect 12139 948 12152 957
rect 12204 948 12217 957
rect 12269 948 12282 957
rect 12334 948 12347 957
rect 11876 914 11909 948
rect 11943 914 11981 948
rect 12015 914 12022 948
rect 12334 914 12341 948
rect 11876 908 12022 914
rect 11876 905 11882 908
rect 12016 905 12022 908
rect 12074 905 12087 914
rect 12139 905 12152 914
rect 12204 905 12217 914
rect 12269 905 12282 914
rect 12334 905 12347 914
rect 12399 905 12412 957
rect 12464 905 12477 957
rect 12529 905 12542 957
rect 12594 905 12607 957
rect 12659 905 12672 957
rect 12724 905 12737 957
rect 12789 905 12802 957
rect 12854 948 12867 957
rect 12919 948 12932 957
rect 12984 948 12997 957
rect 13049 948 13062 957
rect 13114 948 13127 957
rect 13179 948 13192 957
rect 12861 914 12867 948
rect 13114 914 13115 948
rect 13179 914 13187 948
rect 12854 905 12867 914
rect 12919 905 12932 914
rect 12984 905 12997 914
rect 13049 905 13062 914
rect 13114 905 13127 914
rect 13179 905 13192 914
rect 13244 905 13257 957
rect 13309 905 13322 957
rect 13374 905 13387 957
rect 13439 905 13452 957
rect 13504 948 13517 957
rect 13569 948 13582 957
rect 13634 948 13647 957
rect 13699 948 13712 957
rect 13764 948 13777 957
rect 13829 948 13842 957
rect 13509 914 13517 948
rect 13581 914 13582 948
rect 13829 914 13835 948
rect 13504 905 13517 914
rect 13569 905 13582 914
rect 13634 905 13647 914
rect 13699 905 13712 914
rect 13764 905 13777 914
rect 13829 905 13842 914
rect 13894 905 13907 957
rect 13959 905 13972 957
rect 14024 905 14037 957
rect 14089 905 14102 957
rect 14154 948 14167 957
rect 14219 948 14232 957
rect 14284 948 14297 957
rect 14349 948 14362 957
rect 14414 948 14427 957
rect 14479 948 14492 957
rect 14544 948 14557 957
rect 14157 914 14167 948
rect 14229 914 14232 948
rect 14479 914 14483 948
rect 14544 914 14555 948
rect 14154 905 14167 914
rect 14219 905 14232 914
rect 14284 905 14297 914
rect 14349 905 14362 914
rect 14414 905 14427 914
rect 14479 905 14492 914
rect 14544 905 14557 914
rect 14609 905 14622 957
rect 14674 905 14686 957
rect 14738 905 14750 957
rect 14802 948 14814 957
rect 14866 948 14878 957
rect 14930 948 14942 957
rect 14994 948 15006 957
rect 15058 948 15070 957
rect 15122 948 15134 957
rect 14805 914 14814 948
rect 14877 914 14878 948
rect 15058 914 15059 948
rect 15122 914 15131 948
rect 14802 905 14814 914
rect 14866 905 14878 914
rect 14930 905 14942 914
rect 14994 905 15006 914
rect 15058 905 15070 914
rect 15122 905 15134 914
rect 15186 905 15198 957
rect 15250 905 15262 957
rect 15314 905 15326 957
rect 15378 948 15390 957
rect 15442 948 15454 957
rect 15506 948 15518 957
rect 15570 948 15582 957
rect 15634 948 15646 957
rect 15381 914 15390 948
rect 15453 914 15454 948
rect 15634 914 15635 948
rect 15378 905 15390 914
rect 15442 905 15454 914
rect 15506 905 15518 914
rect 15570 905 15582 914
rect 15634 905 15646 914
rect 15698 905 15710 957
rect 15762 905 15774 957
rect 15826 948 15838 957
rect 15826 914 15833 948
rect 15826 905 15838 914
rect 15890 905 15902 957
rect 15954 905 15966 957
rect 16018 905 16030 957
rect 16082 948 16094 957
rect 16146 948 16158 957
rect 16210 948 16222 957
rect 16274 948 16286 957
rect 16338 948 16350 957
rect 16402 948 16414 957
rect 16083 914 16094 948
rect 16155 914 16158 948
rect 16402 914 16409 948
rect 16082 905 16094 914
rect 16146 905 16158 914
rect 16210 905 16222 914
rect 16274 905 16286 914
rect 16338 905 16350 914
rect 16402 905 16414 914
rect 16466 905 16478 957
rect 16530 905 16542 957
rect 16594 905 16606 957
rect 16658 948 16670 957
rect 16722 948 16734 957
rect 16786 948 16798 957
rect 16850 948 16862 957
rect 16914 948 16926 957
rect 16978 948 16990 957
rect 16659 914 16670 948
rect 16731 914 16734 948
rect 16978 914 16985 948
rect 16658 905 16670 914
rect 16722 905 16734 914
rect 16786 905 16798 914
rect 16850 905 16862 914
rect 16914 905 16926 914
rect 16978 905 16990 914
rect 17042 905 17054 957
rect 17106 905 17118 957
rect 17170 905 17182 957
rect 17234 948 17246 957
rect 17298 948 17310 957
rect 17362 948 17374 957
rect 17426 948 17438 957
rect 17490 948 17502 957
rect 17554 948 17566 957
rect 17235 914 17246 948
rect 17307 914 17310 948
rect 17554 914 17561 948
rect 17234 905 17246 914
rect 17298 905 17310 914
rect 17362 905 17374 914
rect 17426 905 17438 914
rect 17490 905 17502 914
rect 17554 905 17566 914
rect 17618 905 17630 957
rect 17682 905 17694 957
rect 17746 905 17758 957
rect 17810 948 17822 957
rect 17874 948 17886 957
rect 17938 948 17950 957
rect 18002 948 18014 957
rect 18066 948 18078 957
rect 18130 948 18142 957
rect 17811 914 17822 948
rect 17883 914 17886 948
rect 18130 914 18137 948
rect 17810 905 17822 914
rect 17874 905 17886 914
rect 17938 905 17950 914
rect 18002 905 18014 914
rect 18066 905 18078 914
rect 18130 905 18142 914
rect 18194 905 18206 957
rect 18258 905 18270 957
rect 18322 905 18334 957
rect 18386 948 18398 957
rect 18450 948 18462 957
rect 18514 948 18526 957
rect 18578 948 18590 957
rect 18642 948 18654 957
rect 18706 948 18718 957
rect 18387 914 18398 948
rect 18459 914 18462 948
rect 18706 914 18713 948
rect 18386 905 18398 914
rect 18450 905 18462 914
rect 18514 905 18526 914
rect 18578 905 18590 914
rect 18642 905 18654 914
rect 18706 905 18718 914
rect 18770 905 18782 957
rect 18834 905 18846 957
rect 18898 905 18910 957
rect 18962 905 18974 957
rect 19026 905 19038 957
rect 19090 905 19102 957
rect 19154 948 19166 957
rect 19218 948 19230 957
rect 19282 948 19294 957
rect 19346 948 19358 957
rect 19410 948 19422 957
rect 19161 914 19166 948
rect 19410 914 19415 948
rect 19154 905 19166 914
rect 19218 905 19230 914
rect 19282 905 19294 914
rect 19346 905 19358 914
rect 19410 905 19422 914
rect 19474 905 19486 957
rect 19538 905 19550 957
rect 19602 905 19614 957
rect 19666 905 19678 957
rect 19730 948 19742 957
rect 19794 948 19806 957
rect 19858 948 19870 957
rect 19922 948 19934 957
rect 19986 948 19998 957
rect 19737 914 19742 948
rect 19986 914 19991 948
rect 19730 905 19742 914
rect 19794 905 19806 914
rect 19858 905 19870 914
rect 19922 905 19934 914
rect 19986 905 19998 914
rect 20050 905 20062 957
rect 20114 905 20126 957
rect 20178 905 20190 957
rect 20242 905 20254 957
rect 20306 948 20318 957
rect 20370 948 20382 957
rect 20434 948 20446 957
rect 20498 948 20510 957
rect 20562 948 20574 957
rect 20313 914 20318 948
rect 20562 914 20567 948
rect 20306 905 20318 914
rect 20370 905 20382 914
rect 20434 905 20446 914
rect 20498 905 20510 914
rect 20562 905 20574 914
rect 20626 905 20638 957
rect 20690 905 20702 957
rect 20754 905 20766 957
rect 20818 905 20830 957
rect 20882 948 20894 957
rect 20946 948 20958 957
rect 21010 948 21022 957
rect 21074 948 21086 957
rect 21138 948 21150 957
rect 20889 914 20894 948
rect 21138 914 21143 948
rect 20882 905 20894 914
rect 20946 905 20958 914
rect 21010 905 21022 914
rect 21074 905 21086 914
rect 21138 905 21150 914
rect 21202 905 21214 957
rect 21266 905 21278 957
rect 21330 905 21342 957
rect 21394 905 21406 957
rect 21458 948 21470 957
rect 21522 948 21534 957
rect 21586 948 21598 957
rect 21650 948 21662 957
rect 21714 948 21726 957
rect 21465 914 21470 948
rect 21714 914 21719 948
rect 21458 905 21470 914
rect 21522 905 21534 914
rect 21586 905 21598 914
rect 21650 905 21662 914
rect 21714 905 21726 914
rect 21778 905 21790 957
rect 21842 905 21854 957
rect 21906 905 21918 957
rect 21970 954 21978 957
tri 21978 954 21981 957 sw
rect 21970 908 21981 954
rect 21970 905 21978 908
tri 21978 905 21981 908 nw
rect 22236 912 22288 915
tri 6313 878 6339 904 sw
rect 22236 902 22248 912
rect 22282 902 22288 912
rect 6267 877 6339 878
tri 6339 877 6340 878 sw
rect 6267 843 6273 877
rect 6307 871 22236 877
rect 6307 843 9388 871
rect 6267 837 9388 843
rect 9422 837 9460 871
rect 9494 837 12538 871
rect 12572 837 12610 871
rect 12644 837 15688 871
rect 15722 837 15760 871
rect 15794 837 18838 871
rect 18872 837 18910 871
rect 18944 837 21988 871
rect 22022 837 22060 871
rect 22094 850 22236 871
rect 22433 864 22439 867
rect 22094 837 22288 850
rect 6267 831 22236 837
rect 1539 824 1545 827
rect 71 818 1545 824
rect 1597 818 1610 827
rect 1662 818 1675 827
rect 1727 818 1740 827
rect 71 784 83 818
rect 117 784 155 818
rect 189 784 227 818
rect 261 784 299 818
rect 333 784 371 818
rect 405 784 443 818
rect 477 784 515 818
rect 549 784 587 818
rect 621 784 659 818
rect 693 784 731 818
rect 765 784 803 818
rect 837 784 875 818
rect 909 784 947 818
rect 981 784 1019 818
rect 1053 784 1091 818
rect 1125 784 1163 818
rect 1197 784 1235 818
rect 1269 784 1307 818
rect 1341 784 1379 818
rect 1413 784 1451 818
rect 1485 784 1523 818
rect 1662 784 1667 818
rect 1727 784 1739 818
rect 71 778 1545 784
rect 1539 775 1545 778
rect 1597 775 1610 784
rect 1662 775 1675 784
rect 1727 775 1740 784
rect 1792 775 1805 827
rect 1857 775 1870 827
rect 1922 775 1935 827
rect 1987 818 2000 827
rect 2052 818 2065 827
rect 2117 818 2130 827
rect 2182 818 2195 827
rect 2247 818 2260 827
rect 2312 818 2325 827
rect 2377 818 2390 827
rect 1989 784 2000 818
rect 2061 784 2065 818
rect 2312 784 2315 818
rect 2377 784 2387 818
rect 1987 775 2000 784
rect 2052 775 2065 784
rect 2117 775 2130 784
rect 2182 775 2195 784
rect 2247 775 2260 784
rect 2312 775 2325 784
rect 2377 775 2390 784
rect 2442 775 2455 827
rect 2507 775 2520 827
rect 2572 775 2585 827
rect 2637 775 2650 827
rect 2702 818 2715 827
rect 2767 818 2780 827
rect 2832 818 2845 827
rect 2897 818 2910 827
rect 2962 818 2975 827
rect 3027 818 3040 827
rect 2709 784 2715 818
rect 2962 784 2963 818
rect 3027 784 3035 818
rect 2702 775 2715 784
rect 2767 775 2780 784
rect 2832 775 2845 784
rect 2897 775 2910 784
rect 2962 775 2975 784
rect 3027 775 3040 784
rect 3092 775 3105 827
rect 3157 775 3170 827
rect 3222 818 3235 827
rect 3222 784 3233 818
rect 3222 775 3235 784
rect 3287 775 3300 827
rect 3352 775 3365 827
rect 3417 775 3430 827
rect 3482 818 3495 827
rect 3547 818 3560 827
rect 3612 818 3625 827
rect 3677 818 3690 827
rect 3742 818 3755 827
rect 3807 818 3820 827
rect 3872 818 3885 827
rect 3483 784 3495 818
rect 3555 784 3560 818
rect 3807 784 3809 818
rect 3872 784 3881 818
rect 3482 775 3495 784
rect 3547 775 3560 784
rect 3612 775 3625 784
rect 3677 775 3690 784
rect 3742 775 3755 784
rect 3807 775 3820 784
rect 3872 775 3885 784
rect 3937 775 3950 827
rect 4002 775 4015 827
rect 4067 775 4080 827
rect 4132 775 4144 827
rect 4196 818 4208 827
rect 4260 818 4272 827
rect 4324 818 4336 827
rect 4388 818 4400 827
rect 4452 818 4464 827
rect 4203 784 4208 818
rect 4452 784 4457 818
rect 4196 775 4208 784
rect 4260 775 4272 784
rect 4324 775 4336 784
rect 4388 775 4400 784
rect 4452 775 4464 784
rect 4516 775 4528 827
rect 4580 775 4592 827
rect 4644 775 4656 827
rect 4708 775 4720 827
rect 4772 818 4784 827
rect 4836 818 4848 827
rect 4900 818 4912 827
rect 4964 818 4976 827
rect 5028 818 5040 827
rect 4779 784 4784 818
rect 5028 784 5033 818
rect 4772 775 4784 784
rect 4836 775 4848 784
rect 4900 775 4912 784
rect 4964 775 4976 784
rect 5028 775 5040 784
rect 5092 775 5104 827
rect 5156 775 5168 827
rect 5220 775 5232 827
rect 5284 775 5296 827
rect 5348 818 5360 827
rect 5412 818 5424 827
rect 5476 818 5488 827
rect 5540 818 5552 827
rect 5604 818 5616 827
rect 5355 784 5360 818
rect 5604 784 5609 818
rect 5348 775 5360 784
rect 5412 775 5424 784
rect 5476 775 5488 784
rect 5540 775 5552 784
rect 5604 775 5616 784
rect 5668 775 5680 827
rect 5732 775 5744 827
rect 5796 775 5808 827
rect 5860 775 5872 827
rect 5924 818 5936 827
rect 5988 818 6000 827
rect 6052 818 6064 827
rect 6116 824 6122 827
rect 6116 818 6231 824
rect 5931 784 5936 818
rect 6147 784 6185 818
rect 6219 784 6231 818
rect 5924 775 5936 784
rect 5988 775 6000 784
rect 6052 775 6064 784
rect 6116 778 6231 784
rect 6267 801 6313 831
tri 6313 804 6340 831 nw
rect 22354 858 22439 864
rect 22354 824 22366 858
rect 22400 824 22438 858
rect 22354 818 22439 824
rect 22433 815 22439 818
rect 22491 815 22507 867
rect 22559 815 22575 867
rect 22627 815 22643 867
rect 22695 815 22711 867
rect 22763 815 22779 867
rect 22831 858 22847 867
rect 22899 858 22915 867
rect 22967 858 22982 867
rect 23034 858 23049 867
rect 23101 858 23116 867
rect 23168 858 23183 867
rect 23235 858 23250 867
rect 23302 864 23308 867
rect 23302 858 24356 864
rect 22832 824 22847 858
rect 22904 824 22915 858
rect 22976 824 22982 858
rect 23048 824 23049 858
rect 23336 824 23374 858
rect 23408 824 23446 858
rect 23480 824 23518 858
rect 23552 824 23590 858
rect 23624 824 23662 858
rect 23696 824 23734 858
rect 23768 824 23806 858
rect 23840 824 23878 858
rect 23912 824 23950 858
rect 23984 824 24022 858
rect 24056 824 24094 858
rect 24128 824 24166 858
rect 24200 824 24238 858
rect 24272 824 24310 858
rect 24344 824 24356 858
rect 22831 815 22847 824
rect 22899 815 22915 824
rect 22967 815 22982 824
rect 23034 815 23049 824
rect 23101 815 23116 824
rect 23168 815 23183 824
rect 23235 815 23250 824
rect 23302 818 24356 824
rect 23302 815 23308 818
rect 6116 775 6122 778
tri 6260 767 6267 774 se
rect 6267 767 6273 801
rect 6307 767 6313 801
rect 7610 798 7616 801
tri 6251 758 6260 767 se
rect 6260 758 6313 767
tri 6240 747 6251 758 se
rect 6251 747 6313 758
rect 6371 792 7616 798
rect 7668 792 7681 801
rect 6371 758 6383 792
rect 6417 758 6455 792
rect 6489 758 6527 792
rect 6561 758 6599 792
rect 6633 758 6671 792
rect 6705 758 6743 792
rect 6777 758 6815 792
rect 6849 758 6887 792
rect 6921 758 6959 792
rect 6993 758 7031 792
rect 7065 758 7103 792
rect 7137 758 7175 792
rect 7209 758 7247 792
rect 7281 758 7319 792
rect 7353 758 7391 792
rect 7425 758 7463 792
rect 7497 758 7535 792
rect 7569 758 7607 792
rect 7668 758 7679 792
rect 6371 752 7616 758
rect 7610 749 7616 752
rect 7668 749 7681 758
rect 7733 749 7746 801
rect 7798 749 7811 801
rect 7863 749 7876 801
rect 7928 792 7941 801
rect 7993 792 8006 801
rect 8058 792 8071 801
rect 8123 792 8136 801
rect 8188 792 8201 801
rect 8253 792 8266 801
rect 8318 792 8331 801
rect 7929 758 7941 792
rect 8001 758 8006 792
rect 8253 758 8255 792
rect 8318 758 8327 792
rect 7928 749 7941 758
rect 7993 749 8006 758
rect 8058 749 8071 758
rect 8123 749 8136 758
rect 8188 749 8201 758
rect 8253 749 8266 758
rect 8318 749 8331 758
rect 8383 749 8396 801
rect 8448 749 8461 801
rect 8513 749 8526 801
rect 8578 749 8591 801
rect 8643 792 8656 801
rect 8708 792 8721 801
rect 8773 792 8786 801
rect 8838 792 8851 801
rect 8903 792 8916 801
rect 8968 792 8981 801
rect 8649 758 8656 792
rect 8968 758 8975 792
rect 8643 749 8656 758
rect 8708 749 8721 758
rect 8773 749 8786 758
rect 8838 749 8851 758
rect 8903 749 8916 758
rect 8968 749 8981 758
rect 9033 749 9046 801
rect 9098 749 9111 801
rect 9163 749 9176 801
rect 9228 749 9241 801
rect 9293 792 9306 801
rect 9358 792 9371 801
rect 9297 758 9306 792
rect 9369 758 9371 792
rect 9293 749 9306 758
rect 9358 749 9371 758
rect 9423 749 9436 801
rect 9488 749 9501 801
rect 9553 792 9566 801
rect 9618 792 9631 801
rect 9683 792 9696 801
rect 9748 792 9761 801
rect 9813 792 9826 801
rect 9748 758 9749 792
rect 9813 758 9821 792
rect 9553 749 9566 758
rect 9618 749 9631 758
rect 9683 749 9696 758
rect 9748 749 9761 758
rect 9813 749 9826 758
rect 9878 749 9891 801
rect 9943 749 9956 801
rect 10008 749 10021 801
rect 10073 749 10086 801
rect 10138 792 10151 801
rect 10203 792 10216 801
rect 10268 792 10281 801
rect 10333 792 10346 801
rect 10398 792 10411 801
rect 10463 792 10476 801
rect 10143 758 10151 792
rect 10215 758 10216 792
rect 10463 758 10469 792
rect 10138 749 10151 758
rect 10203 749 10216 758
rect 10268 749 10281 758
rect 10333 749 10346 758
rect 10398 749 10411 758
rect 10463 749 10476 758
rect 10528 749 10541 801
rect 10593 749 10606 801
rect 10658 749 10671 801
rect 10723 749 10736 801
rect 10788 792 10800 801
rect 10852 792 10864 801
rect 10916 792 10928 801
rect 10980 792 10992 801
rect 11044 792 11056 801
rect 11108 792 11120 801
rect 10791 758 10800 792
rect 10863 758 10864 792
rect 11044 758 11045 792
rect 11108 758 11117 792
rect 10788 749 10800 758
rect 10852 749 10864 758
rect 10916 749 10928 758
rect 10980 749 10992 758
rect 11044 749 11056 758
rect 11108 749 11120 758
rect 11172 749 11184 801
rect 11236 749 11248 801
rect 11300 749 11312 801
rect 11364 792 11376 801
rect 11428 792 11440 801
rect 11492 792 11504 801
rect 11556 792 11568 801
rect 11620 792 11632 801
rect 11684 792 11696 801
rect 11367 758 11376 792
rect 11439 758 11440 792
rect 11620 758 11621 792
rect 11684 758 11693 792
rect 11364 749 11376 758
rect 11428 749 11440 758
rect 11492 749 11504 758
rect 11556 749 11568 758
rect 11620 749 11632 758
rect 11684 749 11696 758
rect 11748 749 11760 801
rect 11812 749 11824 801
rect 11876 798 11882 801
rect 12016 798 12022 801
rect 11876 792 12022 798
rect 12074 792 12087 801
rect 12139 792 12152 801
rect 12204 792 12217 801
rect 12269 792 12282 801
rect 12334 792 12347 801
rect 11876 758 11909 792
rect 11943 758 11981 792
rect 12015 758 12022 792
rect 12334 758 12341 792
rect 11876 752 12022 758
rect 11876 749 11882 752
rect 12016 749 12022 752
rect 12074 749 12087 758
rect 12139 749 12152 758
rect 12204 749 12217 758
rect 12269 749 12282 758
rect 12334 749 12347 758
rect 12399 749 12412 801
rect 12464 749 12477 801
rect 12529 749 12542 801
rect 12594 749 12607 801
rect 12659 749 12672 801
rect 12724 749 12737 801
rect 12789 749 12802 801
rect 12854 792 12867 801
rect 12919 792 12932 801
rect 12984 792 12997 801
rect 13049 792 13062 801
rect 13114 792 13127 801
rect 13179 792 13192 801
rect 12861 758 12867 792
rect 13114 758 13115 792
rect 13179 758 13187 792
rect 12854 749 12867 758
rect 12919 749 12932 758
rect 12984 749 12997 758
rect 13049 749 13062 758
rect 13114 749 13127 758
rect 13179 749 13192 758
rect 13244 749 13257 801
rect 13309 749 13322 801
rect 13374 749 13387 801
rect 13439 749 13452 801
rect 13504 792 13517 801
rect 13569 792 13582 801
rect 13634 792 13647 801
rect 13699 792 13712 801
rect 13764 792 13777 801
rect 13829 792 13842 801
rect 13509 758 13517 792
rect 13581 758 13582 792
rect 13829 758 13835 792
rect 13504 749 13517 758
rect 13569 749 13582 758
rect 13634 749 13647 758
rect 13699 749 13712 758
rect 13764 749 13777 758
rect 13829 749 13842 758
rect 13894 749 13907 801
rect 13959 749 13972 801
rect 14024 749 14037 801
rect 14089 749 14101 801
rect 14153 792 14165 801
rect 14217 792 14229 801
rect 14281 792 14293 801
rect 14345 792 14357 801
rect 14409 792 14421 801
rect 14473 792 14485 801
rect 14157 758 14165 792
rect 14409 758 14411 792
rect 14473 758 14483 792
rect 14153 749 14165 758
rect 14217 749 14229 758
rect 14281 749 14293 758
rect 14345 749 14357 758
rect 14409 749 14421 758
rect 14473 749 14485 758
rect 14537 749 14549 801
rect 14601 749 14613 801
rect 14665 749 14677 801
rect 14729 792 14741 801
rect 14793 792 14805 801
rect 14857 792 14869 801
rect 14921 792 14933 801
rect 14985 792 14997 801
rect 15049 792 15061 801
rect 14733 758 14741 792
rect 14985 758 14987 792
rect 15049 758 15059 792
rect 14729 749 14741 758
rect 14793 749 14805 758
rect 14857 749 14869 758
rect 14921 749 14933 758
rect 14985 749 14997 758
rect 15049 749 15061 758
rect 15113 749 15125 801
rect 15177 749 15189 801
rect 15241 749 15253 801
rect 15305 792 15317 801
rect 15369 792 15381 801
rect 15433 792 15445 801
rect 15497 792 15509 801
rect 15561 792 15573 801
rect 15625 792 15637 801
rect 15309 758 15317 792
rect 15561 758 15563 792
rect 15625 758 15635 792
rect 15305 749 15317 758
rect 15369 749 15381 758
rect 15433 749 15445 758
rect 15497 749 15509 758
rect 15561 749 15573 758
rect 15625 749 15637 758
rect 15689 749 15701 801
rect 15753 749 15765 801
rect 15817 749 15829 801
rect 15881 749 15893 801
rect 15945 749 15957 801
rect 16009 792 16021 801
rect 16073 792 16085 801
rect 16137 792 16149 801
rect 16201 792 16213 801
rect 16265 792 16277 801
rect 16329 792 16341 801
rect 16011 758 16021 792
rect 16083 758 16085 792
rect 16329 758 16337 792
rect 16009 749 16021 758
rect 16073 749 16085 758
rect 16137 749 16149 758
rect 16201 749 16213 758
rect 16265 749 16277 758
rect 16329 749 16341 758
rect 16393 749 16405 801
rect 16457 749 16469 801
rect 16521 749 16533 801
rect 16585 792 16597 801
rect 16649 792 16661 801
rect 16713 792 16725 801
rect 16777 792 16789 801
rect 16841 792 16853 801
rect 16905 792 16917 801
rect 16587 758 16597 792
rect 16659 758 16661 792
rect 16905 758 16913 792
rect 16585 749 16597 758
rect 16649 749 16661 758
rect 16713 749 16725 758
rect 16777 749 16789 758
rect 16841 749 16853 758
rect 16905 749 16917 758
rect 16969 749 16981 801
rect 17033 749 17045 801
rect 17097 749 17109 801
rect 17161 792 17173 801
rect 17225 792 17237 801
rect 17289 792 17301 801
rect 17353 792 17365 801
rect 17417 792 17429 801
rect 17481 792 17493 801
rect 17163 758 17173 792
rect 17235 758 17237 792
rect 17481 758 17489 792
rect 17161 749 17173 758
rect 17225 749 17237 758
rect 17289 749 17301 758
rect 17353 749 17365 758
rect 17417 749 17429 758
rect 17481 749 17493 758
rect 17545 749 17557 801
rect 17609 749 17621 801
rect 17673 749 17685 801
rect 17737 792 17749 801
rect 17801 792 17813 801
rect 17865 792 17877 801
rect 17929 792 17941 801
rect 17993 792 18005 801
rect 18057 792 18069 801
rect 17739 758 17749 792
rect 17811 758 17813 792
rect 18057 758 18065 792
rect 17737 749 17749 758
rect 17801 749 17813 758
rect 17865 749 17877 758
rect 17929 749 17941 758
rect 17993 749 18005 758
rect 18057 749 18069 758
rect 18121 749 18133 801
rect 18185 749 18197 801
rect 18249 749 18261 801
rect 18313 792 18325 801
rect 18377 792 18389 801
rect 18441 792 18453 801
rect 18505 792 18517 801
rect 18569 792 18581 801
rect 18633 792 18645 801
rect 18315 758 18325 792
rect 18387 758 18389 792
rect 18633 758 18641 792
rect 18313 749 18325 758
rect 18377 749 18389 758
rect 18441 749 18453 758
rect 18505 749 18517 758
rect 18569 749 18581 758
rect 18633 749 18645 758
rect 18697 749 18709 801
rect 18761 749 18773 801
rect 18825 749 18837 801
rect 18889 749 18901 801
rect 18953 749 18965 801
rect 19017 749 19029 801
rect 19081 792 19093 801
rect 19145 792 19157 801
rect 19209 792 19221 801
rect 19273 792 19285 801
rect 19337 792 19349 801
rect 19089 758 19093 792
rect 19337 758 19343 792
rect 19081 749 19093 758
rect 19145 749 19157 758
rect 19209 749 19221 758
rect 19273 749 19285 758
rect 19337 749 19349 758
rect 19401 749 19413 801
rect 19465 749 19477 801
rect 19529 749 19541 801
rect 19593 749 19605 801
rect 19657 792 19669 801
rect 19721 792 19733 801
rect 19785 792 19797 801
rect 19849 792 19861 801
rect 19913 792 19925 801
rect 19665 758 19669 792
rect 19913 758 19919 792
rect 19657 749 19669 758
rect 19721 749 19733 758
rect 19785 749 19797 758
rect 19849 749 19861 758
rect 19913 749 19925 758
rect 19977 749 19989 801
rect 20041 749 20053 801
rect 20105 749 20117 801
rect 20169 749 20181 801
rect 20233 792 20245 801
rect 20297 792 20309 801
rect 20361 792 20373 801
rect 20425 792 20437 801
rect 20489 792 20501 801
rect 20241 758 20245 792
rect 20489 758 20495 792
rect 20233 749 20245 758
rect 20297 749 20309 758
rect 20361 749 20373 758
rect 20425 749 20437 758
rect 20489 749 20501 758
rect 20553 749 20565 801
rect 20617 749 20629 801
rect 20681 749 20693 801
rect 20745 749 20757 801
rect 20809 792 20821 801
rect 20873 792 20885 801
rect 20937 792 20949 801
rect 21001 792 21013 801
rect 21065 792 21077 801
rect 20817 758 20821 792
rect 21065 758 21071 792
rect 20809 749 20821 758
rect 20873 749 20885 758
rect 20937 749 20949 758
rect 21001 749 21013 758
rect 21065 749 21077 758
rect 21129 749 21141 801
rect 21193 749 21205 801
rect 21257 749 21269 801
rect 21321 749 21333 801
rect 21385 792 21397 801
rect 21449 792 21461 801
rect 21513 792 21525 801
rect 21577 792 21589 801
rect 21641 792 21653 801
rect 21393 758 21397 792
rect 21641 758 21647 792
rect 21385 749 21397 758
rect 21449 749 21461 758
rect 21513 749 21525 758
rect 21577 749 21589 758
rect 21641 749 21653 758
rect 21705 749 21717 801
rect 21769 749 21781 801
rect 21833 749 21845 801
rect 21897 749 21909 801
rect 21961 798 21967 801
rect 21961 792 21981 798
rect 21969 758 21981 792
rect 21961 752 21981 758
rect 22236 772 22288 785
rect 21961 749 21967 752
rect 72 741 6313 747
rect 72 707 3088 741
rect 3122 707 3160 741
rect 3194 726 6313 741
tri 6313 726 6335 748 sw
rect 3194 725 6335 726
rect 3194 707 6273 725
rect 72 701 6273 707
tri 6245 691 6255 701 ne
rect 6255 691 6273 701
rect 6307 721 6335 725
tri 6335 721 6340 726 sw
rect 6307 720 22236 721
rect 6307 715 22288 720
rect 6307 691 9388 715
tri 6255 681 6265 691 ne
rect 6265 681 9388 691
rect 9422 681 9460 715
rect 9494 681 12538 715
rect 12572 681 12610 715
rect 12644 681 15688 715
rect 15722 681 15760 715
rect 15794 681 18838 715
rect 18872 681 18910 715
rect 18944 681 21988 715
rect 22022 681 22060 715
rect 22094 681 22288 715
tri 23398 708 23401 711 se
rect 23401 708 23407 711
tri 6265 679 6267 681 ne
rect 6267 679 22288 681
tri 6267 675 6271 679 ne
rect 6271 675 22288 679
rect 22354 702 23407 708
rect 23459 702 23478 711
rect 23530 702 23549 711
rect 23601 702 23620 711
rect 23672 702 23691 711
rect 23743 702 23762 711
rect 23814 702 23833 711
rect 23885 702 23904 711
rect 23956 702 23975 711
rect 24027 702 24046 711
rect 24098 708 24104 711
tri 24104 708 24107 711 sw
rect 24098 702 24356 708
rect 1539 668 1545 671
rect 71 662 1545 668
rect 1597 662 1610 671
rect 1662 662 1675 671
rect 1727 662 1740 671
rect 71 628 83 662
rect 117 628 155 662
rect 189 628 227 662
rect 261 628 299 662
rect 333 628 371 662
rect 405 628 443 662
rect 477 628 515 662
rect 549 628 587 662
rect 621 628 659 662
rect 693 628 731 662
rect 765 628 803 662
rect 837 628 875 662
rect 909 628 947 662
rect 981 628 1019 662
rect 1053 628 1091 662
rect 1125 628 1163 662
rect 1197 628 1235 662
rect 1269 628 1307 662
rect 1341 628 1379 662
rect 1413 628 1451 662
rect 1485 628 1523 662
rect 1662 628 1667 662
rect 1727 628 1739 662
rect 71 622 1545 628
rect 1539 619 1545 622
rect 1597 619 1610 628
rect 1662 619 1675 628
rect 1727 619 1740 628
rect 1792 619 1805 671
rect 1857 619 1870 671
rect 1922 619 1935 671
rect 1987 662 2000 671
rect 2052 662 2065 671
rect 2117 662 2130 671
rect 2182 662 2195 671
rect 2247 662 2260 671
rect 2312 662 2325 671
rect 2377 662 2390 671
rect 1989 628 2000 662
rect 2061 628 2065 662
rect 2312 628 2315 662
rect 2377 628 2387 662
rect 1987 619 2000 628
rect 2052 619 2065 628
rect 2117 619 2130 628
rect 2182 619 2195 628
rect 2247 619 2260 628
rect 2312 619 2325 628
rect 2377 619 2390 628
rect 2442 619 2455 671
rect 2507 619 2520 671
rect 2572 619 2585 671
rect 2637 619 2650 671
rect 2702 662 2715 671
rect 2767 662 2780 671
rect 2832 662 2845 671
rect 2897 662 2910 671
rect 2962 662 2975 671
rect 3027 662 3040 671
rect 2709 628 2715 662
rect 2962 628 2963 662
rect 3027 628 3035 662
rect 2702 619 2715 628
rect 2767 619 2780 628
rect 2832 619 2845 628
rect 2897 619 2910 628
rect 2962 619 2975 628
rect 3027 619 3040 628
rect 3092 619 3105 671
rect 3157 619 3170 671
rect 3222 662 3235 671
rect 3222 628 3233 662
rect 3222 619 3235 628
rect 3287 619 3300 671
rect 3352 619 3365 671
rect 3417 619 3430 671
rect 3482 662 3495 671
rect 3547 662 3560 671
rect 3612 662 3625 671
rect 3677 662 3690 671
rect 3742 662 3755 671
rect 3807 662 3820 671
rect 3872 662 3885 671
rect 3483 628 3495 662
rect 3555 628 3560 662
rect 3807 628 3809 662
rect 3872 628 3881 662
rect 3482 619 3495 628
rect 3547 619 3560 628
rect 3612 619 3625 628
rect 3677 619 3690 628
rect 3742 619 3755 628
rect 3807 619 3820 628
rect 3872 619 3885 628
rect 3937 619 3950 671
rect 4002 619 4015 671
rect 4067 619 4080 671
rect 4132 619 4144 671
rect 4196 662 4208 671
rect 4260 662 4272 671
rect 4324 662 4336 671
rect 4388 662 4400 671
rect 4452 662 4464 671
rect 4203 628 4208 662
rect 4452 628 4457 662
rect 4196 619 4208 628
rect 4260 619 4272 628
rect 4324 619 4336 628
rect 4388 619 4400 628
rect 4452 619 4464 628
rect 4516 619 4528 671
rect 4580 619 4592 671
rect 4644 619 4656 671
rect 4708 619 4720 671
rect 4772 662 4784 671
rect 4836 662 4848 671
rect 4900 662 4912 671
rect 4964 662 4976 671
rect 5028 662 5040 671
rect 4779 628 4784 662
rect 5028 628 5033 662
rect 4772 619 4784 628
rect 4836 619 4848 628
rect 4900 619 4912 628
rect 4964 619 4976 628
rect 5028 619 5040 628
rect 5092 619 5104 671
rect 5156 619 5168 671
rect 5220 619 5232 671
rect 5284 619 5296 671
rect 5348 662 5360 671
rect 5412 662 5424 671
rect 5476 662 5488 671
rect 5540 662 5552 671
rect 5604 662 5616 671
rect 5355 628 5360 662
rect 5604 628 5609 662
rect 5348 619 5360 628
rect 5412 619 5424 628
rect 5476 619 5488 628
rect 5540 619 5552 628
rect 5604 619 5616 628
rect 5668 619 5680 671
rect 5732 619 5744 671
rect 5796 619 5808 671
rect 5860 619 5872 671
rect 5924 662 5936 671
rect 5988 662 6000 671
rect 6052 662 6064 671
rect 6116 668 6122 671
rect 22354 668 22366 702
rect 22400 668 22438 702
rect 22472 668 22510 702
rect 22544 668 22582 702
rect 22616 668 22654 702
rect 22688 668 22726 702
rect 22760 668 22798 702
rect 22832 668 22870 702
rect 22904 668 22942 702
rect 22976 668 23014 702
rect 23048 668 23086 702
rect 23120 668 23158 702
rect 23192 668 23230 702
rect 23264 668 23302 702
rect 23336 668 23374 702
rect 24128 668 24166 702
rect 24200 668 24238 702
rect 24272 668 24310 702
rect 24344 668 24356 702
rect 6116 662 6231 668
rect 22354 662 23407 668
rect 5931 628 5936 662
rect 6147 628 6185 662
rect 6219 628 6231 662
tri 23398 659 23401 662 ne
rect 23401 659 23407 662
rect 23459 659 23478 668
rect 23530 659 23549 668
rect 23601 659 23620 668
rect 23672 659 23691 668
rect 23743 659 23762 668
rect 23814 659 23833 668
rect 23885 659 23904 668
rect 23956 659 23975 668
rect 24027 659 24046 668
rect 24098 662 24356 668
rect 24098 659 24104 662
tri 24104 659 24107 662 nw
rect 7610 642 7616 645
rect 5924 619 5936 628
rect 5988 619 6000 628
rect 6052 619 6064 628
rect 6116 622 6231 628
rect 6371 636 7616 642
rect 7668 636 7681 645
rect 6116 619 6122 622
rect 6371 602 6383 636
rect 6417 602 6455 636
rect 6489 602 6527 636
rect 6561 602 6599 636
rect 6633 602 6671 636
rect 6705 602 6743 636
rect 6777 602 6815 636
rect 6849 602 6887 636
rect 6921 602 6959 636
rect 6993 602 7031 636
rect 7065 602 7103 636
rect 7137 602 7175 636
rect 7209 602 7247 636
rect 7281 602 7319 636
rect 7353 602 7391 636
rect 7425 602 7463 636
rect 7497 602 7535 636
rect 7569 602 7607 636
rect 7668 602 7679 636
rect 6371 596 7616 602
rect 7610 593 7616 596
rect 7668 593 7681 602
rect 7733 593 7746 645
rect 7798 593 7811 645
rect 7863 593 7876 645
rect 7928 636 7941 645
rect 7993 636 8006 645
rect 8058 636 8071 645
rect 8123 636 8136 645
rect 8188 636 8201 645
rect 8253 636 8266 645
rect 8318 636 8331 645
rect 7929 602 7941 636
rect 8001 602 8006 636
rect 8253 602 8255 636
rect 8318 602 8327 636
rect 7928 593 7941 602
rect 7993 593 8006 602
rect 8058 593 8071 602
rect 8123 593 8136 602
rect 8188 593 8201 602
rect 8253 593 8266 602
rect 8318 593 8331 602
rect 8383 593 8396 645
rect 8448 593 8461 645
rect 8513 593 8526 645
rect 8578 593 8591 645
rect 8643 636 8656 645
rect 8708 636 8721 645
rect 8773 636 8786 645
rect 8838 636 8851 645
rect 8903 636 8916 645
rect 8968 636 8981 645
rect 8649 602 8656 636
rect 8968 602 8975 636
rect 8643 593 8656 602
rect 8708 593 8721 602
rect 8773 593 8786 602
rect 8838 593 8851 602
rect 8903 593 8916 602
rect 8968 593 8981 602
rect 9033 593 9046 645
rect 9098 593 9111 645
rect 9163 593 9176 645
rect 9228 593 9241 645
rect 9293 636 9306 645
rect 9358 636 9371 645
rect 9297 602 9306 636
rect 9369 602 9371 636
rect 9293 593 9306 602
rect 9358 593 9371 602
rect 9423 593 9436 645
rect 9488 593 9501 645
rect 9553 636 9566 645
rect 9618 636 9631 645
rect 9683 636 9696 645
rect 9748 636 9761 645
rect 9813 636 9826 645
rect 9748 602 9749 636
rect 9813 602 9821 636
rect 9553 593 9566 602
rect 9618 593 9631 602
rect 9683 593 9696 602
rect 9748 593 9761 602
rect 9813 593 9826 602
rect 9878 593 9891 645
rect 9943 593 9956 645
rect 10008 593 10021 645
rect 10073 593 10086 645
rect 10138 636 10151 645
rect 10203 636 10216 645
rect 10268 636 10281 645
rect 10333 636 10346 645
rect 10398 636 10411 645
rect 10463 636 10476 645
rect 10143 602 10151 636
rect 10215 602 10216 636
rect 10463 602 10469 636
rect 10138 593 10151 602
rect 10203 593 10216 602
rect 10268 593 10281 602
rect 10333 593 10346 602
rect 10398 593 10411 602
rect 10463 593 10476 602
rect 10528 593 10541 645
rect 10593 593 10606 645
rect 10658 593 10671 645
rect 10723 593 10736 645
rect 10788 636 10800 645
rect 10852 636 10864 645
rect 10916 636 10928 645
rect 10980 636 10992 645
rect 11044 636 11056 645
rect 11108 636 11120 645
rect 10791 602 10800 636
rect 10863 602 10864 636
rect 11044 602 11045 636
rect 11108 602 11117 636
rect 10788 593 10800 602
rect 10852 593 10864 602
rect 10916 593 10928 602
rect 10980 593 10992 602
rect 11044 593 11056 602
rect 11108 593 11120 602
rect 11172 593 11184 645
rect 11236 593 11248 645
rect 11300 593 11312 645
rect 11364 636 11376 645
rect 11428 636 11440 645
rect 11492 636 11504 645
rect 11556 636 11568 645
rect 11620 636 11632 645
rect 11684 636 11696 645
rect 11367 602 11376 636
rect 11439 602 11440 636
rect 11620 602 11621 636
rect 11684 602 11693 636
rect 11364 593 11376 602
rect 11428 593 11440 602
rect 11492 593 11504 602
rect 11556 593 11568 602
rect 11620 593 11632 602
rect 11684 593 11696 602
rect 11748 593 11760 645
rect 11812 593 11824 645
rect 11876 642 11882 645
rect 12016 642 12022 645
rect 11876 636 12022 642
rect 12074 636 12087 645
rect 12139 636 12152 645
rect 12204 636 12217 645
rect 12269 636 12282 645
rect 12334 636 12347 645
rect 11876 602 11909 636
rect 11943 602 11981 636
rect 12015 602 12022 636
rect 12334 602 12341 636
rect 11876 596 12022 602
rect 11876 593 11882 596
rect 12016 593 12022 596
rect 12074 593 12087 602
rect 12139 593 12152 602
rect 12204 593 12217 602
rect 12269 593 12282 602
rect 12334 593 12347 602
rect 12399 593 12412 645
rect 12464 593 12477 645
rect 12529 593 12542 645
rect 12594 593 12607 645
rect 12659 593 12672 645
rect 12724 593 12737 645
rect 12789 593 12802 645
rect 12854 636 12867 645
rect 12919 636 12932 645
rect 12984 636 12997 645
rect 13049 636 13062 645
rect 13114 636 13127 645
rect 13179 636 13192 645
rect 12861 602 12867 636
rect 13114 602 13115 636
rect 13179 602 13187 636
rect 12854 593 12867 602
rect 12919 593 12932 602
rect 12984 593 12997 602
rect 13049 593 13062 602
rect 13114 593 13127 602
rect 13179 593 13192 602
rect 13244 593 13257 645
rect 13309 593 13322 645
rect 13374 593 13387 645
rect 13439 593 13452 645
rect 13504 636 13517 645
rect 13569 636 13582 645
rect 13634 636 13647 645
rect 13699 636 13712 645
rect 13764 636 13777 645
rect 13829 636 13842 645
rect 13509 602 13517 636
rect 13581 602 13582 636
rect 13829 602 13835 636
rect 13504 593 13517 602
rect 13569 593 13582 602
rect 13634 593 13647 602
rect 13699 593 13712 602
rect 13764 593 13777 602
rect 13829 593 13842 602
rect 13894 593 13907 645
rect 13959 593 13972 645
rect 14024 593 14037 645
rect 14089 593 14102 645
rect 14154 636 14167 645
rect 14219 636 14232 645
rect 14284 636 14297 645
rect 14349 636 14362 645
rect 14414 636 14427 645
rect 14479 636 14492 645
rect 14544 636 14557 645
rect 14157 602 14167 636
rect 14229 602 14232 636
rect 14479 602 14483 636
rect 14544 602 14555 636
rect 14154 593 14167 602
rect 14219 593 14232 602
rect 14284 593 14297 602
rect 14349 593 14362 602
rect 14414 593 14427 602
rect 14479 593 14492 602
rect 14544 593 14557 602
rect 14609 593 14622 645
rect 14674 593 14687 645
rect 14739 593 14752 645
rect 14804 636 14817 645
rect 14869 636 14882 645
rect 14934 636 14947 645
rect 14999 636 15012 645
rect 15064 636 15077 645
rect 15129 636 15142 645
rect 15194 636 15206 645
rect 14805 602 14817 636
rect 14877 602 14882 636
rect 15129 602 15131 636
rect 15194 602 15203 636
rect 14804 593 14817 602
rect 14869 593 14882 602
rect 14934 593 14947 602
rect 14999 593 15012 602
rect 15064 593 15077 602
rect 15129 593 15142 602
rect 15194 593 15206 602
rect 15258 593 15270 645
rect 15322 593 15334 645
rect 15386 593 15398 645
rect 15450 636 15462 645
rect 15514 636 15526 645
rect 15578 636 15590 645
rect 15642 636 15654 645
rect 15453 602 15462 636
rect 15525 602 15526 636
rect 15450 593 15462 602
rect 15514 593 15526 602
rect 15578 593 15590 602
rect 15642 593 15654 602
rect 15706 593 15718 645
rect 15770 593 15782 645
rect 15834 636 15846 645
rect 15898 636 15910 645
rect 15898 602 15905 636
rect 15834 593 15846 602
rect 15898 593 15910 602
rect 15962 593 15974 645
rect 16026 593 16038 645
rect 16090 593 16102 645
rect 16154 636 16166 645
rect 16218 636 16230 645
rect 16282 636 16294 645
rect 16346 636 16358 645
rect 16410 636 16422 645
rect 16474 636 16486 645
rect 16155 602 16166 636
rect 16227 602 16230 636
rect 16474 602 16481 636
rect 16154 593 16166 602
rect 16218 593 16230 602
rect 16282 593 16294 602
rect 16346 593 16358 602
rect 16410 593 16422 602
rect 16474 593 16486 602
rect 16538 593 16550 645
rect 16602 593 16614 645
rect 16666 593 16678 645
rect 16730 636 16742 645
rect 16794 636 16806 645
rect 16858 636 16870 645
rect 16922 636 16934 645
rect 16986 636 16998 645
rect 17050 636 17062 645
rect 16731 602 16742 636
rect 16803 602 16806 636
rect 17050 602 17057 636
rect 16730 593 16742 602
rect 16794 593 16806 602
rect 16858 593 16870 602
rect 16922 593 16934 602
rect 16986 593 16998 602
rect 17050 593 17062 602
rect 17114 593 17126 645
rect 17178 593 17190 645
rect 17242 593 17254 645
rect 17306 636 17318 645
rect 17370 636 17382 645
rect 17434 636 17446 645
rect 17498 636 17510 645
rect 17562 636 17574 645
rect 17626 636 17638 645
rect 17307 602 17318 636
rect 17379 602 17382 636
rect 17626 602 17633 636
rect 17306 593 17318 602
rect 17370 593 17382 602
rect 17434 593 17446 602
rect 17498 593 17510 602
rect 17562 593 17574 602
rect 17626 593 17638 602
rect 17690 593 17702 645
rect 17754 593 17766 645
rect 17818 593 17830 645
rect 17882 636 17894 645
rect 17946 636 17958 645
rect 18010 636 18022 645
rect 18074 636 18086 645
rect 18138 636 18150 645
rect 18202 636 18214 645
rect 17883 602 17894 636
rect 17955 602 17958 636
rect 18202 602 18209 636
rect 17882 593 17894 602
rect 17946 593 17958 602
rect 18010 593 18022 602
rect 18074 593 18086 602
rect 18138 593 18150 602
rect 18202 593 18214 602
rect 18266 593 18278 645
rect 18330 593 18342 645
rect 18394 593 18406 645
rect 18458 636 18470 645
rect 18522 636 18534 645
rect 18586 636 18598 645
rect 18650 636 18662 645
rect 18714 636 18726 645
rect 18778 636 18790 645
rect 18459 602 18470 636
rect 18531 602 18534 636
rect 18778 602 18785 636
rect 18458 593 18470 602
rect 18522 593 18534 602
rect 18586 593 18598 602
rect 18650 593 18662 602
rect 18714 593 18726 602
rect 18778 593 18790 602
rect 18842 593 18854 645
rect 18906 593 18918 645
rect 18970 593 18982 645
rect 19034 593 19046 645
rect 19098 593 19110 645
rect 19162 593 19174 645
rect 19226 636 19238 645
rect 19290 636 19302 645
rect 19354 636 19366 645
rect 19418 636 19430 645
rect 19482 636 19494 645
rect 19233 602 19238 636
rect 19482 602 19487 636
rect 19226 593 19238 602
rect 19290 593 19302 602
rect 19354 593 19366 602
rect 19418 593 19430 602
rect 19482 593 19494 602
rect 19546 593 19558 645
rect 19610 593 19622 645
rect 19674 593 19686 645
rect 19738 593 19750 645
rect 19802 636 19814 645
rect 19866 636 19878 645
rect 19930 636 19942 645
rect 19994 636 20006 645
rect 20058 636 20070 645
rect 19809 602 19814 636
rect 20058 602 20063 636
rect 19802 593 19814 602
rect 19866 593 19878 602
rect 19930 593 19942 602
rect 19994 593 20006 602
rect 20058 593 20070 602
rect 20122 593 20134 645
rect 20186 593 20198 645
rect 20250 593 20262 645
rect 20314 593 20326 645
rect 20378 636 20390 645
rect 20442 636 20454 645
rect 20506 636 20518 645
rect 20570 636 20582 645
rect 20634 636 20646 645
rect 20385 602 20390 636
rect 20634 602 20639 636
rect 20378 593 20390 602
rect 20442 593 20454 602
rect 20506 593 20518 602
rect 20570 593 20582 602
rect 20634 593 20646 602
rect 20698 593 20710 645
rect 20762 593 20774 645
rect 20826 593 20838 645
rect 20890 593 20902 645
rect 20954 636 20966 645
rect 21018 636 21030 645
rect 21082 636 21094 645
rect 21146 636 21158 645
rect 21210 636 21222 645
rect 20961 602 20966 636
rect 21210 602 21215 636
rect 20954 593 20966 602
rect 21018 593 21030 602
rect 21082 593 21094 602
rect 21146 593 21158 602
rect 21210 593 21222 602
rect 21274 593 21286 645
rect 21338 593 21350 645
rect 21402 593 21414 645
rect 21466 593 21478 645
rect 21530 636 21542 645
rect 21594 636 21606 645
rect 21658 636 21670 645
rect 21722 636 21734 645
rect 21786 636 21798 645
rect 21537 602 21542 636
rect 21786 602 21791 636
rect 21530 593 21542 602
rect 21594 593 21606 602
rect 21658 593 21670 602
rect 21722 593 21734 602
rect 21786 593 21798 602
rect 21850 593 21862 645
rect 21914 593 21926 645
rect 21978 593 21984 645
rect 20688 473 20694 525
rect 20746 473 20760 525
rect 20812 473 20826 525
rect 20878 473 20892 525
rect 20944 473 20957 525
rect 21009 473 21022 525
rect 21074 473 21080 525
rect 20688 461 21080 473
rect 20688 409 20694 461
rect 20746 409 20760 461
rect 20812 409 20826 461
rect 20878 409 20892 461
rect 20944 409 20957 461
rect 21009 409 21022 461
rect 21074 409 21080 461
rect 20688 397 21080 409
rect 20688 345 20694 397
rect 20746 345 20760 397
rect 20812 345 20826 397
rect 20878 345 20892 397
rect 20944 345 20957 397
rect 21009 345 21022 397
rect 21074 345 21080 397
rect 23401 473 23407 525
rect 23459 473 23478 525
rect 23530 473 23549 525
rect 23601 473 23620 525
rect 23672 473 23691 525
rect 23743 473 23761 525
rect 23813 473 23831 525
rect 23883 473 23901 525
rect 23953 473 23971 525
rect 24023 473 24041 525
rect 24093 473 24099 525
rect 23401 461 24099 473
rect 23401 409 23407 461
rect 23459 409 23478 461
rect 23530 409 23549 461
rect 23601 409 23620 461
rect 23672 409 23691 461
rect 23743 409 23761 461
rect 23813 409 23831 461
rect 23883 409 23901 461
rect 23953 409 23971 461
rect 24023 409 24041 461
rect 24093 409 24099 461
rect 23401 397 24099 409
rect 23401 345 23407 397
rect 23459 345 23478 397
rect 23530 345 23549 397
rect 23601 345 23620 397
rect 23672 345 23691 397
rect 23743 345 23761 397
rect 23813 345 23831 397
rect 23883 345 23901 397
rect 23953 345 23971 397
rect 24023 345 24041 397
rect 24093 345 24099 397
<< via1 >>
rect 22436 2106 22488 2115
rect 22436 2072 22438 2106
rect 22438 2072 22472 2106
rect 22472 2072 22488 2106
rect 22436 2063 22488 2072
rect 22504 2106 22556 2115
rect 22504 2072 22510 2106
rect 22510 2072 22544 2106
rect 22544 2072 22556 2106
rect 22504 2063 22556 2072
rect 22572 2106 22624 2115
rect 22572 2072 22582 2106
rect 22582 2072 22616 2106
rect 22616 2072 22624 2106
rect 22572 2063 22624 2072
rect 22640 2106 22692 2115
rect 22640 2072 22654 2106
rect 22654 2072 22688 2106
rect 22688 2072 22692 2106
rect 22640 2063 22692 2072
rect 22708 2106 22760 2115
rect 22708 2072 22726 2106
rect 22726 2072 22760 2106
rect 22708 2063 22760 2072
rect 22776 2106 22828 2115
rect 22844 2106 22896 2115
rect 22912 2106 22964 2115
rect 22980 2106 23032 2115
rect 23048 2106 23100 2115
rect 23116 2106 23168 2115
rect 23183 2106 23235 2115
rect 23250 2106 23302 2115
rect 22776 2072 22798 2106
rect 22798 2072 22828 2106
rect 22844 2072 22870 2106
rect 22870 2072 22896 2106
rect 22912 2072 22942 2106
rect 22942 2072 22964 2106
rect 22980 2072 23014 2106
rect 23014 2072 23032 2106
rect 23048 2072 23086 2106
rect 23086 2072 23100 2106
rect 23116 2072 23120 2106
rect 23120 2072 23158 2106
rect 23158 2072 23168 2106
rect 23183 2072 23192 2106
rect 23192 2072 23230 2106
rect 23230 2072 23235 2106
rect 23250 2072 23264 2106
rect 23264 2072 23302 2106
rect 22776 2063 22828 2072
rect 22844 2063 22896 2072
rect 22912 2063 22964 2072
rect 22980 2063 23032 2072
rect 23048 2063 23100 2072
rect 23116 2063 23168 2072
rect 23183 2063 23235 2072
rect 23250 2063 23302 2072
rect 22236 2049 22288 2055
rect 22236 2015 22248 2049
rect 22248 2015 22282 2049
rect 22282 2015 22288 2049
rect 22236 2003 22288 2015
rect 22236 1974 22288 1991
rect 22236 1940 22248 1974
rect 22248 1940 22282 1974
rect 22282 1940 22288 1974
rect 22236 1939 22288 1940
rect 22236 1899 22288 1927
rect 23407 1950 23459 1959
rect 23478 1950 23530 1959
rect 23549 1950 23601 1959
rect 23620 1950 23672 1959
rect 23691 1950 23743 1959
rect 23762 1950 23814 1959
rect 23833 1950 23885 1959
rect 23904 1950 23956 1959
rect 23975 1950 24027 1959
rect 24046 1950 24098 1959
rect 23407 1916 23408 1950
rect 23408 1916 23446 1950
rect 23446 1916 23459 1950
rect 23478 1916 23480 1950
rect 23480 1916 23518 1950
rect 23518 1916 23530 1950
rect 23549 1916 23552 1950
rect 23552 1916 23590 1950
rect 23590 1916 23601 1950
rect 23620 1916 23624 1950
rect 23624 1916 23662 1950
rect 23662 1916 23672 1950
rect 23691 1916 23696 1950
rect 23696 1916 23734 1950
rect 23734 1916 23743 1950
rect 23762 1916 23768 1950
rect 23768 1916 23806 1950
rect 23806 1916 23814 1950
rect 23833 1916 23840 1950
rect 23840 1916 23878 1950
rect 23878 1916 23885 1950
rect 23904 1916 23912 1950
rect 23912 1916 23950 1950
rect 23950 1916 23956 1950
rect 23975 1916 23984 1950
rect 23984 1916 24022 1950
rect 24022 1916 24027 1950
rect 24046 1916 24056 1950
rect 24056 1916 24094 1950
rect 24094 1916 24098 1950
rect 23407 1907 23459 1916
rect 23478 1907 23530 1916
rect 23549 1907 23601 1916
rect 23620 1907 23672 1916
rect 23691 1907 23743 1916
rect 23762 1907 23814 1916
rect 23833 1907 23885 1916
rect 23904 1907 23956 1916
rect 23975 1907 24027 1916
rect 24046 1907 24098 1916
rect 22236 1875 22248 1899
rect 22248 1875 22282 1899
rect 22282 1875 22288 1899
rect 22236 1824 22288 1863
rect 22236 1811 22248 1824
rect 22248 1811 22282 1824
rect 22282 1811 22288 1824
rect 22236 1790 22248 1799
rect 22248 1790 22282 1799
rect 22282 1790 22288 1799
rect 22236 1748 22288 1790
rect 22439 1794 22491 1803
rect 22439 1760 22472 1794
rect 22472 1760 22491 1794
rect 22439 1751 22491 1760
rect 22507 1794 22559 1803
rect 22507 1760 22510 1794
rect 22510 1760 22544 1794
rect 22544 1760 22559 1794
rect 22507 1751 22559 1760
rect 22575 1794 22627 1803
rect 22575 1760 22582 1794
rect 22582 1760 22616 1794
rect 22616 1760 22627 1794
rect 22575 1751 22627 1760
rect 22643 1794 22695 1803
rect 22643 1760 22654 1794
rect 22654 1760 22688 1794
rect 22688 1760 22695 1794
rect 22643 1751 22695 1760
rect 22711 1794 22763 1803
rect 22711 1760 22726 1794
rect 22726 1760 22760 1794
rect 22760 1760 22763 1794
rect 22711 1751 22763 1760
rect 22779 1794 22831 1803
rect 22847 1794 22899 1803
rect 22915 1794 22967 1803
rect 22982 1794 23034 1803
rect 23049 1794 23101 1803
rect 23116 1794 23168 1803
rect 23183 1794 23235 1803
rect 23250 1794 23302 1803
rect 22779 1760 22798 1794
rect 22798 1760 22831 1794
rect 22847 1760 22870 1794
rect 22870 1760 22899 1794
rect 22915 1760 22942 1794
rect 22942 1760 22967 1794
rect 22982 1760 23014 1794
rect 23014 1760 23034 1794
rect 23049 1760 23086 1794
rect 23086 1760 23101 1794
rect 23116 1760 23120 1794
rect 23120 1760 23158 1794
rect 23158 1760 23168 1794
rect 23183 1760 23192 1794
rect 23192 1760 23230 1794
rect 23230 1760 23235 1794
rect 23250 1760 23264 1794
rect 23264 1760 23302 1794
rect 22779 1751 22831 1760
rect 22847 1751 22899 1760
rect 22915 1751 22967 1760
rect 22982 1751 23034 1760
rect 23049 1751 23101 1760
rect 23116 1751 23168 1760
rect 23183 1751 23235 1760
rect 23250 1751 23302 1760
rect 22236 1747 22248 1748
rect 22248 1747 22282 1748
rect 22282 1747 22288 1748
rect 22236 1714 22248 1735
rect 22248 1714 22282 1735
rect 22282 1714 22288 1735
rect 22236 1683 22288 1714
rect 22236 1638 22248 1671
rect 22248 1638 22282 1671
rect 22282 1638 22288 1671
rect 22236 1619 22288 1638
rect 22236 1596 22288 1607
rect 23407 1638 23459 1647
rect 23478 1638 23530 1647
rect 23549 1638 23601 1647
rect 23620 1638 23672 1647
rect 23691 1638 23743 1647
rect 23762 1638 23814 1647
rect 23833 1638 23885 1647
rect 23904 1638 23956 1647
rect 23975 1638 24027 1647
rect 24046 1638 24098 1647
rect 23407 1604 23408 1638
rect 23408 1604 23446 1638
rect 23446 1604 23459 1638
rect 23478 1604 23480 1638
rect 23480 1604 23518 1638
rect 23518 1604 23530 1638
rect 23549 1604 23552 1638
rect 23552 1604 23590 1638
rect 23590 1604 23601 1638
rect 23620 1604 23624 1638
rect 23624 1604 23662 1638
rect 23662 1604 23672 1638
rect 23691 1604 23696 1638
rect 23696 1604 23734 1638
rect 23734 1604 23743 1638
rect 23762 1604 23768 1638
rect 23768 1604 23806 1638
rect 23806 1604 23814 1638
rect 23833 1604 23840 1638
rect 23840 1604 23878 1638
rect 23878 1604 23885 1638
rect 23904 1604 23912 1638
rect 23912 1604 23950 1638
rect 23950 1604 23956 1638
rect 23975 1604 23984 1638
rect 23984 1604 24022 1638
rect 24022 1604 24027 1638
rect 24046 1604 24056 1638
rect 24056 1604 24094 1638
rect 24094 1604 24098 1638
rect 22236 1562 22248 1596
rect 22248 1562 22282 1596
rect 22282 1562 22288 1596
rect 23407 1595 23459 1604
rect 23478 1595 23530 1604
rect 23549 1595 23601 1604
rect 23620 1595 23672 1604
rect 23691 1595 23743 1604
rect 23762 1595 23814 1604
rect 23833 1595 23885 1604
rect 23904 1595 23956 1604
rect 23975 1595 24027 1604
rect 24046 1595 24098 1604
rect 22236 1555 22288 1562
rect 22236 1520 22288 1543
rect 22236 1491 22248 1520
rect 22248 1491 22282 1520
rect 22282 1491 22288 1520
rect 22236 1444 22288 1479
rect 22236 1427 22248 1444
rect 22248 1427 22282 1444
rect 22282 1427 22288 1444
rect 22439 1482 22491 1491
rect 22439 1448 22472 1482
rect 22472 1448 22491 1482
rect 22439 1439 22491 1448
rect 22507 1482 22559 1491
rect 22507 1448 22510 1482
rect 22510 1448 22544 1482
rect 22544 1448 22559 1482
rect 22507 1439 22559 1448
rect 22575 1482 22627 1491
rect 22575 1448 22582 1482
rect 22582 1448 22616 1482
rect 22616 1448 22627 1482
rect 22575 1439 22627 1448
rect 22643 1482 22695 1491
rect 22643 1448 22654 1482
rect 22654 1448 22688 1482
rect 22688 1448 22695 1482
rect 22643 1439 22695 1448
rect 22711 1482 22763 1491
rect 22711 1448 22726 1482
rect 22726 1448 22760 1482
rect 22760 1448 22763 1482
rect 22711 1439 22763 1448
rect 22779 1482 22831 1491
rect 22847 1482 22899 1491
rect 22915 1482 22967 1491
rect 22982 1482 23034 1491
rect 23049 1482 23101 1491
rect 23116 1482 23168 1491
rect 23183 1482 23235 1491
rect 23250 1482 23302 1491
rect 22779 1448 22798 1482
rect 22798 1448 22831 1482
rect 22847 1448 22870 1482
rect 22870 1448 22899 1482
rect 22915 1448 22942 1482
rect 22942 1448 22967 1482
rect 22982 1448 23014 1482
rect 23014 1448 23034 1482
rect 23049 1448 23086 1482
rect 23086 1448 23101 1482
rect 23116 1448 23120 1482
rect 23120 1448 23158 1482
rect 23158 1448 23168 1482
rect 23183 1448 23192 1482
rect 23192 1448 23230 1482
rect 23230 1448 23235 1482
rect 23250 1448 23264 1482
rect 23264 1448 23302 1482
rect 22779 1439 22831 1448
rect 22847 1439 22899 1448
rect 22915 1439 22967 1448
rect 22982 1439 23034 1448
rect 23049 1439 23101 1448
rect 23116 1439 23168 1448
rect 23183 1439 23235 1448
rect 23250 1439 23302 1448
rect 22236 1410 22248 1415
rect 22248 1410 22282 1415
rect 22282 1410 22288 1415
rect 22236 1368 22288 1410
rect 22236 1363 22248 1368
rect 22248 1363 22282 1368
rect 22282 1363 22288 1368
rect 22236 1334 22248 1351
rect 22248 1334 22282 1351
rect 22282 1334 22288 1351
rect 22236 1299 22288 1334
rect 7616 1260 7668 1269
rect 7681 1260 7733 1269
rect 7616 1226 7641 1260
rect 7641 1226 7668 1260
rect 7681 1226 7713 1260
rect 7713 1226 7733 1260
rect 7616 1217 7668 1226
rect 7681 1217 7733 1226
rect 7746 1260 7798 1269
rect 7746 1226 7751 1260
rect 7751 1226 7785 1260
rect 7785 1226 7798 1260
rect 7746 1217 7798 1226
rect 7811 1260 7863 1269
rect 7811 1226 7823 1260
rect 7823 1226 7857 1260
rect 7857 1226 7863 1260
rect 7811 1217 7863 1226
rect 7876 1260 7928 1269
rect 7941 1260 7993 1269
rect 8006 1260 8058 1269
rect 8071 1260 8123 1269
rect 8136 1260 8188 1269
rect 8201 1260 8253 1269
rect 8266 1260 8318 1269
rect 8331 1260 8383 1269
rect 7876 1226 7895 1260
rect 7895 1226 7928 1260
rect 7941 1226 7967 1260
rect 7967 1226 7993 1260
rect 8006 1226 8039 1260
rect 8039 1226 8058 1260
rect 8071 1226 8073 1260
rect 8073 1226 8111 1260
rect 8111 1226 8123 1260
rect 8136 1226 8145 1260
rect 8145 1226 8183 1260
rect 8183 1226 8188 1260
rect 8201 1226 8217 1260
rect 8217 1226 8253 1260
rect 8266 1226 8289 1260
rect 8289 1226 8318 1260
rect 8331 1226 8361 1260
rect 8361 1226 8383 1260
rect 7876 1217 7928 1226
rect 7941 1217 7993 1226
rect 8006 1217 8058 1226
rect 8071 1217 8123 1226
rect 8136 1217 8188 1226
rect 8201 1217 8253 1226
rect 8266 1217 8318 1226
rect 8331 1217 8383 1226
rect 8396 1260 8448 1269
rect 8396 1226 8399 1260
rect 8399 1226 8433 1260
rect 8433 1226 8448 1260
rect 8396 1217 8448 1226
rect 8461 1260 8513 1269
rect 8461 1226 8471 1260
rect 8471 1226 8505 1260
rect 8505 1226 8513 1260
rect 8461 1217 8513 1226
rect 8526 1260 8578 1269
rect 8526 1226 8543 1260
rect 8543 1226 8577 1260
rect 8577 1226 8578 1260
rect 8526 1217 8578 1226
rect 8591 1260 8643 1269
rect 8656 1260 8708 1269
rect 8721 1260 8773 1269
rect 8786 1260 8838 1269
rect 8851 1260 8903 1269
rect 8916 1260 8968 1269
rect 8981 1260 9033 1269
rect 8591 1226 8615 1260
rect 8615 1226 8643 1260
rect 8656 1226 8687 1260
rect 8687 1226 8708 1260
rect 8721 1226 8759 1260
rect 8759 1226 8773 1260
rect 8786 1226 8793 1260
rect 8793 1226 8831 1260
rect 8831 1226 8838 1260
rect 8851 1226 8865 1260
rect 8865 1226 8903 1260
rect 8916 1226 8937 1260
rect 8937 1226 8968 1260
rect 8981 1226 9009 1260
rect 9009 1226 9033 1260
rect 8591 1217 8643 1226
rect 8656 1217 8708 1226
rect 8721 1217 8773 1226
rect 8786 1217 8838 1226
rect 8851 1217 8903 1226
rect 8916 1217 8968 1226
rect 8981 1217 9033 1226
rect 9046 1260 9098 1269
rect 9046 1226 9047 1260
rect 9047 1226 9081 1260
rect 9081 1226 9098 1260
rect 9046 1217 9098 1226
rect 9111 1260 9163 1269
rect 9111 1226 9119 1260
rect 9119 1226 9153 1260
rect 9153 1226 9163 1260
rect 9111 1217 9163 1226
rect 9176 1260 9228 1269
rect 9176 1226 9191 1260
rect 9191 1226 9225 1260
rect 9225 1226 9228 1260
rect 9176 1217 9228 1226
rect 9241 1260 9293 1269
rect 9306 1260 9358 1269
rect 9241 1226 9263 1260
rect 9263 1226 9293 1260
rect 9306 1226 9335 1260
rect 9335 1226 9358 1260
rect 9241 1217 9293 1226
rect 9306 1217 9358 1226
rect 9371 1217 9423 1269
rect 9436 1217 9488 1269
rect 9501 1260 9553 1269
rect 9566 1260 9618 1269
rect 9631 1260 9683 1269
rect 9696 1260 9748 1269
rect 9761 1260 9813 1269
rect 9826 1260 9878 1269
rect 9501 1226 9533 1260
rect 9533 1226 9553 1260
rect 9566 1226 9567 1260
rect 9567 1226 9605 1260
rect 9605 1226 9618 1260
rect 9631 1226 9639 1260
rect 9639 1226 9677 1260
rect 9677 1226 9683 1260
rect 9696 1226 9711 1260
rect 9711 1226 9748 1260
rect 9761 1226 9783 1260
rect 9783 1226 9813 1260
rect 9826 1226 9855 1260
rect 9855 1226 9878 1260
rect 9501 1217 9553 1226
rect 9566 1217 9618 1226
rect 9631 1217 9683 1226
rect 9696 1217 9748 1226
rect 9761 1217 9813 1226
rect 9826 1217 9878 1226
rect 9891 1260 9943 1269
rect 9891 1226 9893 1260
rect 9893 1226 9927 1260
rect 9927 1226 9943 1260
rect 9891 1217 9943 1226
rect 9956 1260 10008 1269
rect 9956 1226 9965 1260
rect 9965 1226 9999 1260
rect 9999 1226 10008 1260
rect 9956 1217 10008 1226
rect 10021 1260 10073 1269
rect 10021 1226 10037 1260
rect 10037 1226 10071 1260
rect 10071 1226 10073 1260
rect 10021 1217 10073 1226
rect 10086 1260 10138 1269
rect 10151 1260 10203 1269
rect 10216 1260 10268 1269
rect 10281 1260 10333 1269
rect 10346 1260 10398 1269
rect 10411 1260 10463 1269
rect 10476 1260 10528 1269
rect 10086 1226 10109 1260
rect 10109 1226 10138 1260
rect 10151 1226 10181 1260
rect 10181 1226 10203 1260
rect 10216 1226 10253 1260
rect 10253 1226 10268 1260
rect 10281 1226 10287 1260
rect 10287 1226 10325 1260
rect 10325 1226 10333 1260
rect 10346 1226 10359 1260
rect 10359 1226 10397 1260
rect 10397 1226 10398 1260
rect 10411 1226 10431 1260
rect 10431 1226 10463 1260
rect 10476 1226 10503 1260
rect 10503 1226 10528 1260
rect 10086 1217 10138 1226
rect 10151 1217 10203 1226
rect 10216 1217 10268 1226
rect 10281 1217 10333 1226
rect 10346 1217 10398 1226
rect 10411 1217 10463 1226
rect 10476 1217 10528 1226
rect 10541 1260 10593 1269
rect 10541 1226 10575 1260
rect 10575 1226 10593 1260
rect 10541 1217 10593 1226
rect 10606 1260 10658 1269
rect 10606 1226 10613 1260
rect 10613 1226 10647 1260
rect 10647 1226 10658 1260
rect 10606 1217 10658 1226
rect 10671 1260 10723 1269
rect 10671 1226 10685 1260
rect 10685 1226 10719 1260
rect 10719 1226 10723 1260
rect 10671 1217 10723 1226
rect 10736 1260 10788 1269
rect 10800 1260 10852 1269
rect 10864 1260 10916 1269
rect 10928 1260 10980 1269
rect 10992 1260 11044 1269
rect 11056 1260 11108 1269
rect 11120 1260 11172 1269
rect 10736 1226 10757 1260
rect 10757 1226 10788 1260
rect 10800 1226 10829 1260
rect 10829 1226 10852 1260
rect 10864 1226 10901 1260
rect 10901 1226 10916 1260
rect 10928 1226 10935 1260
rect 10935 1226 10973 1260
rect 10973 1226 10980 1260
rect 10992 1226 11007 1260
rect 11007 1226 11044 1260
rect 11056 1226 11079 1260
rect 11079 1226 11108 1260
rect 11120 1226 11151 1260
rect 11151 1226 11172 1260
rect 10736 1217 10788 1226
rect 10800 1217 10852 1226
rect 10864 1217 10916 1226
rect 10928 1217 10980 1226
rect 10992 1217 11044 1226
rect 11056 1217 11108 1226
rect 11120 1217 11172 1226
rect 11184 1260 11236 1269
rect 11184 1226 11189 1260
rect 11189 1226 11223 1260
rect 11223 1226 11236 1260
rect 11184 1217 11236 1226
rect 11248 1260 11300 1269
rect 11248 1226 11261 1260
rect 11261 1226 11295 1260
rect 11295 1226 11300 1260
rect 11248 1217 11300 1226
rect 11312 1260 11364 1269
rect 11376 1260 11428 1269
rect 11440 1260 11492 1269
rect 11504 1260 11556 1269
rect 11568 1260 11620 1269
rect 11632 1260 11684 1269
rect 11696 1260 11748 1269
rect 11312 1226 11333 1260
rect 11333 1226 11364 1260
rect 11376 1226 11405 1260
rect 11405 1226 11428 1260
rect 11440 1226 11477 1260
rect 11477 1226 11492 1260
rect 11504 1226 11511 1260
rect 11511 1226 11549 1260
rect 11549 1226 11556 1260
rect 11568 1226 11583 1260
rect 11583 1226 11620 1260
rect 11632 1226 11655 1260
rect 11655 1226 11684 1260
rect 11696 1226 11727 1260
rect 11727 1226 11748 1260
rect 11312 1217 11364 1226
rect 11376 1217 11428 1226
rect 11440 1217 11492 1226
rect 11504 1217 11556 1226
rect 11568 1217 11620 1226
rect 11632 1217 11684 1226
rect 11696 1217 11748 1226
rect 11760 1260 11812 1269
rect 11760 1226 11765 1260
rect 11765 1226 11799 1260
rect 11799 1226 11812 1260
rect 11760 1217 11812 1226
rect 11824 1260 11876 1269
rect 11824 1226 11837 1260
rect 11837 1226 11871 1260
rect 11871 1226 11876 1260
rect 11824 1217 11876 1226
rect 12594 1218 12646 1270
rect 12659 1260 12711 1270
rect 12724 1260 12776 1270
rect 12789 1260 12841 1270
rect 12854 1260 12906 1270
rect 12919 1260 12971 1270
rect 12984 1260 13036 1270
rect 13049 1260 13101 1270
rect 12659 1226 12683 1260
rect 12683 1226 12711 1260
rect 12724 1226 12755 1260
rect 12755 1226 12776 1260
rect 12789 1226 12827 1260
rect 12827 1226 12841 1260
rect 12854 1226 12861 1260
rect 12861 1226 12899 1260
rect 12899 1226 12906 1260
rect 12919 1226 12933 1260
rect 12933 1226 12971 1260
rect 12984 1226 13005 1260
rect 13005 1226 13036 1260
rect 13049 1226 13077 1260
rect 13077 1226 13101 1260
rect 12659 1218 12711 1226
rect 12724 1218 12776 1226
rect 12789 1218 12841 1226
rect 12854 1218 12906 1226
rect 12919 1218 12971 1226
rect 12984 1218 13036 1226
rect 13049 1218 13101 1226
rect 13114 1260 13166 1270
rect 13114 1226 13115 1260
rect 13115 1226 13149 1260
rect 13149 1226 13166 1260
rect 13114 1218 13166 1226
rect 13179 1260 13231 1270
rect 13179 1226 13187 1260
rect 13187 1226 13221 1260
rect 13221 1226 13231 1260
rect 13179 1218 13231 1226
rect 13244 1260 13296 1270
rect 13244 1226 13259 1260
rect 13259 1226 13293 1260
rect 13293 1226 13296 1260
rect 13244 1218 13296 1226
rect 13309 1260 13361 1270
rect 13374 1260 13426 1270
rect 13439 1260 13491 1270
rect 13504 1260 13556 1270
rect 13569 1260 13621 1270
rect 13633 1260 13685 1270
rect 13697 1260 13749 1270
rect 13309 1226 13331 1260
rect 13331 1226 13361 1260
rect 13374 1226 13403 1260
rect 13403 1226 13426 1260
rect 13439 1226 13475 1260
rect 13475 1226 13491 1260
rect 13504 1226 13509 1260
rect 13509 1226 13547 1260
rect 13547 1226 13556 1260
rect 13569 1226 13581 1260
rect 13581 1226 13619 1260
rect 13619 1226 13621 1260
rect 13633 1226 13653 1260
rect 13653 1226 13685 1260
rect 13697 1226 13725 1260
rect 13725 1226 13749 1260
rect 13309 1218 13361 1226
rect 13374 1218 13426 1226
rect 13439 1218 13491 1226
rect 13504 1218 13556 1226
rect 13569 1218 13621 1226
rect 13633 1218 13685 1226
rect 13697 1218 13749 1226
rect 13761 1260 13813 1270
rect 13761 1226 13763 1260
rect 13763 1226 13797 1260
rect 13797 1226 13813 1260
rect 13761 1218 13813 1226
rect 13825 1260 13877 1270
rect 13825 1226 13835 1260
rect 13835 1226 13869 1260
rect 13869 1226 13877 1260
rect 13825 1218 13877 1226
rect 13889 1260 13941 1270
rect 13889 1226 13907 1260
rect 13907 1226 13941 1260
rect 13889 1218 13941 1226
rect 13953 1260 14005 1270
rect 14017 1260 14069 1270
rect 14081 1260 14133 1270
rect 14145 1260 14197 1270
rect 14209 1260 14261 1270
rect 14273 1260 14325 1270
rect 13953 1226 13979 1260
rect 13979 1226 14005 1260
rect 14017 1226 14051 1260
rect 14051 1226 14069 1260
rect 14081 1226 14085 1260
rect 14085 1226 14123 1260
rect 14123 1226 14133 1260
rect 14145 1226 14157 1260
rect 14157 1226 14195 1260
rect 14195 1226 14197 1260
rect 14209 1226 14229 1260
rect 14229 1226 14261 1260
rect 14273 1226 14301 1260
rect 14301 1226 14325 1260
rect 13953 1218 14005 1226
rect 14017 1218 14069 1226
rect 14081 1218 14133 1226
rect 14145 1218 14197 1226
rect 14209 1218 14261 1226
rect 14273 1218 14325 1226
rect 14337 1260 14389 1270
rect 14337 1226 14339 1260
rect 14339 1226 14373 1260
rect 14373 1226 14389 1260
rect 14337 1218 14389 1226
rect 14401 1260 14453 1270
rect 14401 1226 14411 1260
rect 14411 1226 14445 1260
rect 14445 1226 14453 1260
rect 14401 1218 14453 1226
rect 14465 1260 14517 1270
rect 14465 1226 14483 1260
rect 14483 1226 14517 1260
rect 14465 1218 14517 1226
rect 14529 1260 14581 1270
rect 14593 1260 14645 1270
rect 14657 1260 14709 1270
rect 14721 1260 14773 1270
rect 14785 1260 14837 1270
rect 14849 1260 14901 1270
rect 14529 1226 14555 1260
rect 14555 1226 14581 1260
rect 14593 1226 14627 1260
rect 14627 1226 14645 1260
rect 14657 1226 14661 1260
rect 14661 1226 14699 1260
rect 14699 1226 14709 1260
rect 14721 1226 14733 1260
rect 14733 1226 14771 1260
rect 14771 1226 14773 1260
rect 14785 1226 14805 1260
rect 14805 1226 14837 1260
rect 14849 1226 14877 1260
rect 14877 1226 14901 1260
rect 14529 1218 14581 1226
rect 14593 1218 14645 1226
rect 14657 1218 14709 1226
rect 14721 1218 14773 1226
rect 14785 1218 14837 1226
rect 14849 1218 14901 1226
rect 14913 1260 14965 1270
rect 14913 1226 14915 1260
rect 14915 1226 14949 1260
rect 14949 1226 14965 1260
rect 14913 1218 14965 1226
rect 14977 1260 15029 1270
rect 14977 1226 14987 1260
rect 14987 1226 15021 1260
rect 15021 1226 15029 1260
rect 14977 1218 15029 1226
rect 15041 1260 15093 1270
rect 15041 1226 15059 1260
rect 15059 1226 15093 1260
rect 15041 1218 15093 1226
rect 15105 1260 15157 1270
rect 15169 1260 15221 1270
rect 15233 1260 15285 1270
rect 15297 1260 15349 1270
rect 15361 1260 15413 1270
rect 15425 1260 15477 1270
rect 15105 1226 15131 1260
rect 15131 1226 15157 1260
rect 15169 1226 15203 1260
rect 15203 1226 15221 1260
rect 15233 1226 15237 1260
rect 15237 1226 15275 1260
rect 15275 1226 15285 1260
rect 15297 1226 15309 1260
rect 15309 1226 15347 1260
rect 15347 1226 15349 1260
rect 15361 1226 15381 1260
rect 15381 1226 15413 1260
rect 15425 1226 15453 1260
rect 15453 1226 15477 1260
rect 15105 1218 15157 1226
rect 15169 1218 15221 1226
rect 15233 1218 15285 1226
rect 15297 1218 15349 1226
rect 15361 1218 15413 1226
rect 15425 1218 15477 1226
rect 15489 1260 15541 1270
rect 15489 1226 15491 1260
rect 15491 1226 15525 1260
rect 15525 1226 15541 1260
rect 15489 1218 15541 1226
rect 15553 1260 15605 1270
rect 15553 1226 15563 1260
rect 15563 1226 15597 1260
rect 15597 1226 15605 1260
rect 15553 1218 15605 1226
rect 15617 1260 15669 1270
rect 15617 1226 15635 1260
rect 15635 1226 15669 1260
rect 15617 1218 15669 1226
rect 15681 1218 15733 1270
rect 15745 1218 15797 1270
rect 15809 1260 15861 1270
rect 15873 1260 15925 1270
rect 15937 1260 15989 1270
rect 16001 1260 16053 1270
rect 16065 1260 16117 1270
rect 16129 1260 16181 1270
rect 15809 1226 15833 1260
rect 15833 1226 15861 1260
rect 15873 1226 15905 1260
rect 15905 1226 15925 1260
rect 15937 1226 15939 1260
rect 15939 1226 15977 1260
rect 15977 1226 15989 1260
rect 16001 1226 16011 1260
rect 16011 1226 16049 1260
rect 16049 1226 16053 1260
rect 16065 1226 16083 1260
rect 16083 1226 16117 1260
rect 16129 1226 16155 1260
rect 16155 1226 16181 1260
rect 15809 1218 15861 1226
rect 15873 1218 15925 1226
rect 15937 1218 15989 1226
rect 16001 1218 16053 1226
rect 16065 1218 16117 1226
rect 16129 1218 16181 1226
rect 16193 1260 16245 1270
rect 16193 1226 16227 1260
rect 16227 1226 16245 1260
rect 16193 1218 16245 1226
rect 16257 1260 16309 1270
rect 16257 1226 16265 1260
rect 16265 1226 16299 1260
rect 16299 1226 16309 1260
rect 16257 1218 16309 1226
rect 16321 1260 16373 1270
rect 16321 1226 16337 1260
rect 16337 1226 16371 1260
rect 16371 1226 16373 1260
rect 16321 1218 16373 1226
rect 16385 1260 16437 1270
rect 16449 1260 16501 1270
rect 16513 1260 16565 1270
rect 16577 1260 16629 1270
rect 16641 1260 16693 1270
rect 16705 1260 16757 1270
rect 16385 1226 16409 1260
rect 16409 1226 16437 1260
rect 16449 1226 16481 1260
rect 16481 1226 16501 1260
rect 16513 1226 16515 1260
rect 16515 1226 16553 1260
rect 16553 1226 16565 1260
rect 16577 1226 16587 1260
rect 16587 1226 16625 1260
rect 16625 1226 16629 1260
rect 16641 1226 16659 1260
rect 16659 1226 16693 1260
rect 16705 1226 16731 1260
rect 16731 1226 16757 1260
rect 16385 1218 16437 1226
rect 16449 1218 16501 1226
rect 16513 1218 16565 1226
rect 16577 1218 16629 1226
rect 16641 1218 16693 1226
rect 16705 1218 16757 1226
rect 16769 1260 16821 1270
rect 16769 1226 16803 1260
rect 16803 1226 16821 1260
rect 16769 1218 16821 1226
rect 16833 1260 16885 1270
rect 16833 1226 16841 1260
rect 16841 1226 16875 1260
rect 16875 1226 16885 1260
rect 16833 1218 16885 1226
rect 16897 1260 16949 1270
rect 16897 1226 16913 1260
rect 16913 1226 16947 1260
rect 16947 1226 16949 1260
rect 16897 1218 16949 1226
rect 16961 1260 17013 1270
rect 17025 1260 17077 1270
rect 17089 1260 17141 1270
rect 17153 1260 17205 1270
rect 17217 1260 17269 1270
rect 17281 1260 17333 1270
rect 16961 1226 16985 1260
rect 16985 1226 17013 1260
rect 17025 1226 17057 1260
rect 17057 1226 17077 1260
rect 17089 1226 17091 1260
rect 17091 1226 17129 1260
rect 17129 1226 17141 1260
rect 17153 1226 17163 1260
rect 17163 1226 17201 1260
rect 17201 1226 17205 1260
rect 17217 1226 17235 1260
rect 17235 1226 17269 1260
rect 17281 1226 17307 1260
rect 17307 1226 17333 1260
rect 16961 1218 17013 1226
rect 17025 1218 17077 1226
rect 17089 1218 17141 1226
rect 17153 1218 17205 1226
rect 17217 1218 17269 1226
rect 17281 1218 17333 1226
rect 17345 1260 17397 1270
rect 17345 1226 17379 1260
rect 17379 1226 17397 1260
rect 17345 1218 17397 1226
rect 17409 1260 17461 1270
rect 17409 1226 17417 1260
rect 17417 1226 17451 1260
rect 17451 1226 17461 1260
rect 17409 1218 17461 1226
rect 17473 1260 17525 1270
rect 17473 1226 17489 1260
rect 17489 1226 17523 1260
rect 17523 1226 17525 1260
rect 17473 1218 17525 1226
rect 17537 1260 17589 1270
rect 17601 1260 17653 1270
rect 17665 1260 17717 1270
rect 17729 1260 17781 1270
rect 17793 1260 17845 1270
rect 17857 1260 17909 1270
rect 17537 1226 17561 1260
rect 17561 1226 17589 1260
rect 17601 1226 17633 1260
rect 17633 1226 17653 1260
rect 17665 1226 17667 1260
rect 17667 1226 17705 1260
rect 17705 1226 17717 1260
rect 17729 1226 17739 1260
rect 17739 1226 17777 1260
rect 17777 1226 17781 1260
rect 17793 1226 17811 1260
rect 17811 1226 17845 1260
rect 17857 1226 17883 1260
rect 17883 1226 17909 1260
rect 17537 1218 17589 1226
rect 17601 1218 17653 1226
rect 17665 1218 17717 1226
rect 17729 1218 17781 1226
rect 17793 1218 17845 1226
rect 17857 1218 17909 1226
rect 17921 1260 17973 1270
rect 17921 1226 17955 1260
rect 17955 1226 17973 1260
rect 17921 1218 17973 1226
rect 17985 1260 18037 1270
rect 17985 1226 17993 1260
rect 17993 1226 18027 1260
rect 18027 1226 18037 1260
rect 17985 1218 18037 1226
rect 18049 1260 18101 1270
rect 18049 1226 18065 1260
rect 18065 1226 18099 1260
rect 18099 1226 18101 1260
rect 18049 1218 18101 1226
rect 18113 1260 18165 1270
rect 18177 1260 18229 1270
rect 18241 1260 18293 1270
rect 18305 1260 18357 1270
rect 18369 1260 18421 1270
rect 18433 1260 18485 1270
rect 18113 1226 18137 1260
rect 18137 1226 18165 1260
rect 18177 1226 18209 1260
rect 18209 1226 18229 1260
rect 18241 1226 18243 1260
rect 18243 1226 18281 1260
rect 18281 1226 18293 1260
rect 18305 1226 18315 1260
rect 18315 1226 18353 1260
rect 18353 1226 18357 1260
rect 18369 1226 18387 1260
rect 18387 1226 18421 1260
rect 18433 1226 18459 1260
rect 18459 1226 18485 1260
rect 18113 1218 18165 1226
rect 18177 1218 18229 1226
rect 18241 1218 18293 1226
rect 18305 1218 18357 1226
rect 18369 1218 18421 1226
rect 18433 1218 18485 1226
rect 18497 1260 18549 1270
rect 18497 1226 18531 1260
rect 18531 1226 18549 1260
rect 18497 1218 18549 1226
rect 18561 1260 18613 1270
rect 18561 1226 18569 1260
rect 18569 1226 18603 1260
rect 18603 1226 18613 1260
rect 18561 1218 18613 1226
rect 18625 1260 18677 1270
rect 18625 1226 18641 1260
rect 18641 1226 18675 1260
rect 18675 1226 18677 1260
rect 18625 1218 18677 1226
rect 18689 1260 18741 1270
rect 18753 1260 18805 1270
rect 18817 1260 18869 1270
rect 18689 1226 18713 1260
rect 18713 1226 18741 1260
rect 18753 1226 18785 1260
rect 18785 1226 18805 1260
rect 18817 1226 18819 1260
rect 18819 1226 18869 1260
rect 18689 1218 18741 1226
rect 18753 1218 18805 1226
rect 18817 1218 18869 1226
rect 18881 1218 18933 1270
rect 18945 1260 18997 1270
rect 19009 1260 19061 1270
rect 19073 1260 19125 1270
rect 19137 1260 19189 1270
rect 19201 1260 19253 1270
rect 18945 1226 18983 1260
rect 18983 1226 18997 1260
rect 19009 1226 19017 1260
rect 19017 1226 19055 1260
rect 19055 1226 19061 1260
rect 19073 1226 19089 1260
rect 19089 1226 19125 1260
rect 19137 1226 19161 1260
rect 19161 1226 19189 1260
rect 19201 1226 19233 1260
rect 19233 1226 19253 1260
rect 18945 1218 18997 1226
rect 19009 1218 19061 1226
rect 19073 1218 19125 1226
rect 19137 1218 19189 1226
rect 19201 1218 19253 1226
rect 19265 1260 19317 1270
rect 19265 1226 19271 1260
rect 19271 1226 19305 1260
rect 19305 1226 19317 1260
rect 19265 1218 19317 1226
rect 19329 1260 19381 1270
rect 19329 1226 19343 1260
rect 19343 1226 19377 1260
rect 19377 1226 19381 1260
rect 19329 1218 19381 1226
rect 19393 1260 19445 1270
rect 19457 1260 19509 1270
rect 19521 1260 19573 1270
rect 19585 1260 19637 1270
rect 19649 1260 19701 1270
rect 19713 1260 19765 1270
rect 19777 1260 19829 1270
rect 19393 1226 19415 1260
rect 19415 1226 19445 1260
rect 19457 1226 19487 1260
rect 19487 1226 19509 1260
rect 19521 1226 19559 1260
rect 19559 1226 19573 1260
rect 19585 1226 19593 1260
rect 19593 1226 19631 1260
rect 19631 1226 19637 1260
rect 19649 1226 19665 1260
rect 19665 1226 19701 1260
rect 19713 1226 19737 1260
rect 19737 1226 19765 1260
rect 19777 1226 19809 1260
rect 19809 1226 19829 1260
rect 19393 1218 19445 1226
rect 19457 1218 19509 1226
rect 19521 1218 19573 1226
rect 19585 1218 19637 1226
rect 19649 1218 19701 1226
rect 19713 1218 19765 1226
rect 19777 1218 19829 1226
rect 19841 1260 19893 1270
rect 19841 1226 19847 1260
rect 19847 1226 19881 1260
rect 19881 1226 19893 1260
rect 19841 1218 19893 1226
rect 19905 1260 19957 1270
rect 19905 1226 19919 1260
rect 19919 1226 19953 1260
rect 19953 1226 19957 1260
rect 19905 1218 19957 1226
rect 19969 1260 20021 1270
rect 20033 1260 20085 1270
rect 20097 1260 20149 1270
rect 20161 1260 20213 1270
rect 20225 1260 20277 1270
rect 20289 1260 20341 1270
rect 20353 1260 20405 1270
rect 19969 1226 19991 1260
rect 19991 1226 20021 1260
rect 20033 1226 20063 1260
rect 20063 1226 20085 1260
rect 20097 1226 20135 1260
rect 20135 1226 20149 1260
rect 20161 1226 20169 1260
rect 20169 1226 20207 1260
rect 20207 1226 20213 1260
rect 20225 1226 20241 1260
rect 20241 1226 20277 1260
rect 20289 1226 20313 1260
rect 20313 1226 20341 1260
rect 20353 1226 20385 1260
rect 20385 1226 20405 1260
rect 19969 1218 20021 1226
rect 20033 1218 20085 1226
rect 20097 1218 20149 1226
rect 20161 1218 20213 1226
rect 20225 1218 20277 1226
rect 20289 1218 20341 1226
rect 20353 1218 20405 1226
rect 20417 1260 20469 1270
rect 20417 1226 20423 1260
rect 20423 1226 20457 1260
rect 20457 1226 20469 1260
rect 20417 1218 20469 1226
rect 20481 1260 20533 1270
rect 20481 1226 20495 1260
rect 20495 1226 20529 1260
rect 20529 1226 20533 1260
rect 20481 1218 20533 1226
rect 20545 1260 20597 1270
rect 20609 1260 20661 1270
rect 20673 1260 20725 1270
rect 20737 1260 20789 1270
rect 20801 1260 20853 1270
rect 20865 1260 20917 1270
rect 20929 1260 20981 1270
rect 20545 1226 20567 1260
rect 20567 1226 20597 1260
rect 20609 1226 20639 1260
rect 20639 1226 20661 1260
rect 20673 1226 20711 1260
rect 20711 1226 20725 1260
rect 20737 1226 20745 1260
rect 20745 1226 20783 1260
rect 20783 1226 20789 1260
rect 20801 1226 20817 1260
rect 20817 1226 20853 1260
rect 20865 1226 20889 1260
rect 20889 1226 20917 1260
rect 20929 1226 20961 1260
rect 20961 1226 20981 1260
rect 20545 1218 20597 1226
rect 20609 1218 20661 1226
rect 20673 1218 20725 1226
rect 20737 1218 20789 1226
rect 20801 1218 20853 1226
rect 20865 1218 20917 1226
rect 20929 1218 20981 1226
rect 20993 1260 21045 1270
rect 20993 1226 20999 1260
rect 20999 1226 21033 1260
rect 21033 1226 21045 1260
rect 20993 1218 21045 1226
rect 21057 1260 21109 1270
rect 21057 1226 21071 1260
rect 21071 1226 21105 1260
rect 21105 1226 21109 1260
rect 21057 1218 21109 1226
rect 21121 1260 21173 1270
rect 21185 1260 21237 1270
rect 21249 1260 21301 1270
rect 21313 1260 21365 1270
rect 21377 1260 21429 1270
rect 21441 1260 21493 1270
rect 21505 1260 21557 1270
rect 21121 1226 21143 1260
rect 21143 1226 21173 1260
rect 21185 1226 21215 1260
rect 21215 1226 21237 1260
rect 21249 1226 21287 1260
rect 21287 1226 21301 1260
rect 21313 1226 21321 1260
rect 21321 1226 21359 1260
rect 21359 1226 21365 1260
rect 21377 1226 21393 1260
rect 21393 1226 21429 1260
rect 21441 1226 21465 1260
rect 21465 1226 21493 1260
rect 21505 1226 21537 1260
rect 21537 1226 21557 1260
rect 21121 1218 21173 1226
rect 21185 1218 21237 1226
rect 21249 1218 21301 1226
rect 21313 1218 21365 1226
rect 21377 1218 21429 1226
rect 21441 1218 21493 1226
rect 21505 1218 21557 1226
rect 21569 1260 21621 1270
rect 21569 1226 21575 1260
rect 21575 1226 21609 1260
rect 21609 1226 21621 1260
rect 21569 1218 21621 1226
rect 21633 1260 21685 1270
rect 21633 1226 21647 1260
rect 21647 1226 21681 1260
rect 21681 1226 21685 1260
rect 21633 1218 21685 1226
rect 21697 1260 21749 1270
rect 21761 1260 21813 1270
rect 21825 1260 21877 1270
rect 21889 1260 21941 1270
rect 21697 1226 21719 1260
rect 21719 1226 21749 1260
rect 21761 1226 21791 1260
rect 21791 1226 21813 1260
rect 21825 1226 21863 1260
rect 21863 1226 21877 1260
rect 21889 1226 21897 1260
rect 21897 1226 21935 1260
rect 21935 1226 21941 1260
rect 21697 1218 21749 1226
rect 21761 1218 21813 1226
rect 21825 1218 21877 1226
rect 21889 1218 21941 1226
rect 22236 1258 22248 1287
rect 22248 1258 22282 1287
rect 22282 1258 22288 1287
rect 23407 1326 23459 1335
rect 23478 1326 23530 1335
rect 23549 1326 23601 1335
rect 23620 1326 23672 1335
rect 23691 1326 23743 1335
rect 23762 1326 23814 1335
rect 23833 1326 23885 1335
rect 23904 1326 23956 1335
rect 23975 1326 24027 1335
rect 24046 1326 24098 1335
rect 23407 1292 23408 1326
rect 23408 1292 23446 1326
rect 23446 1292 23459 1326
rect 23478 1292 23480 1326
rect 23480 1292 23518 1326
rect 23518 1292 23530 1326
rect 23549 1292 23552 1326
rect 23552 1292 23590 1326
rect 23590 1292 23601 1326
rect 23620 1292 23624 1326
rect 23624 1292 23662 1326
rect 23662 1292 23672 1326
rect 23691 1292 23696 1326
rect 23696 1292 23734 1326
rect 23734 1292 23743 1326
rect 23762 1292 23768 1326
rect 23768 1292 23806 1326
rect 23806 1292 23814 1326
rect 23833 1292 23840 1326
rect 23840 1292 23878 1326
rect 23878 1292 23885 1326
rect 23904 1292 23912 1326
rect 23912 1292 23950 1326
rect 23950 1292 23956 1326
rect 23975 1292 23984 1326
rect 23984 1292 24022 1326
rect 24022 1292 24027 1326
rect 24046 1292 24056 1326
rect 24056 1292 24094 1326
rect 24094 1292 24098 1326
rect 23407 1283 23459 1292
rect 23478 1283 23530 1292
rect 23549 1283 23601 1292
rect 23620 1283 23672 1292
rect 23691 1283 23743 1292
rect 23762 1283 23814 1292
rect 23833 1283 23885 1292
rect 23904 1283 23956 1292
rect 23975 1283 24027 1292
rect 24046 1283 24098 1292
rect 22236 1235 22288 1258
rect 22236 1216 22288 1223
rect 22236 1182 22248 1216
rect 22248 1182 22282 1216
rect 22282 1182 22288 1216
rect 22236 1171 22288 1182
rect 22236 1140 22288 1159
rect 7616 1104 7668 1113
rect 7681 1104 7733 1113
rect 7616 1070 7641 1104
rect 7641 1070 7668 1104
rect 7681 1070 7713 1104
rect 7713 1070 7733 1104
rect 7616 1061 7668 1070
rect 7681 1061 7733 1070
rect 7746 1104 7798 1113
rect 7746 1070 7751 1104
rect 7751 1070 7785 1104
rect 7785 1070 7798 1104
rect 7746 1061 7798 1070
rect 7811 1104 7863 1113
rect 7811 1070 7823 1104
rect 7823 1070 7857 1104
rect 7857 1070 7863 1104
rect 7811 1061 7863 1070
rect 7876 1104 7928 1113
rect 7941 1104 7993 1113
rect 8006 1104 8058 1113
rect 8071 1104 8123 1113
rect 8136 1104 8188 1113
rect 8201 1104 8253 1113
rect 8266 1104 8318 1113
rect 8331 1104 8383 1113
rect 7876 1070 7895 1104
rect 7895 1070 7928 1104
rect 7941 1070 7967 1104
rect 7967 1070 7993 1104
rect 8006 1070 8039 1104
rect 8039 1070 8058 1104
rect 8071 1070 8073 1104
rect 8073 1070 8111 1104
rect 8111 1070 8123 1104
rect 8136 1070 8145 1104
rect 8145 1070 8183 1104
rect 8183 1070 8188 1104
rect 8201 1070 8217 1104
rect 8217 1070 8253 1104
rect 8266 1070 8289 1104
rect 8289 1070 8318 1104
rect 8331 1070 8361 1104
rect 8361 1070 8383 1104
rect 7876 1061 7928 1070
rect 7941 1061 7993 1070
rect 8006 1061 8058 1070
rect 8071 1061 8123 1070
rect 8136 1061 8188 1070
rect 8201 1061 8253 1070
rect 8266 1061 8318 1070
rect 8331 1061 8383 1070
rect 8396 1104 8448 1113
rect 8396 1070 8399 1104
rect 8399 1070 8433 1104
rect 8433 1070 8448 1104
rect 8396 1061 8448 1070
rect 8461 1104 8513 1113
rect 8461 1070 8471 1104
rect 8471 1070 8505 1104
rect 8505 1070 8513 1104
rect 8461 1061 8513 1070
rect 8526 1104 8578 1113
rect 8526 1070 8543 1104
rect 8543 1070 8577 1104
rect 8577 1070 8578 1104
rect 8526 1061 8578 1070
rect 8591 1104 8643 1113
rect 8656 1104 8708 1113
rect 8721 1104 8773 1113
rect 8786 1104 8838 1113
rect 8851 1104 8903 1113
rect 8916 1104 8968 1113
rect 8981 1104 9033 1113
rect 8591 1070 8615 1104
rect 8615 1070 8643 1104
rect 8656 1070 8687 1104
rect 8687 1070 8708 1104
rect 8721 1070 8759 1104
rect 8759 1070 8773 1104
rect 8786 1070 8793 1104
rect 8793 1070 8831 1104
rect 8831 1070 8838 1104
rect 8851 1070 8865 1104
rect 8865 1070 8903 1104
rect 8916 1070 8937 1104
rect 8937 1070 8968 1104
rect 8981 1070 9009 1104
rect 9009 1070 9033 1104
rect 8591 1061 8643 1070
rect 8656 1061 8708 1070
rect 8721 1061 8773 1070
rect 8786 1061 8838 1070
rect 8851 1061 8903 1070
rect 8916 1061 8968 1070
rect 8981 1061 9033 1070
rect 9046 1104 9098 1113
rect 9046 1070 9047 1104
rect 9047 1070 9081 1104
rect 9081 1070 9098 1104
rect 9046 1061 9098 1070
rect 9111 1104 9163 1113
rect 9111 1070 9119 1104
rect 9119 1070 9153 1104
rect 9153 1070 9163 1104
rect 9111 1061 9163 1070
rect 9176 1104 9228 1113
rect 9176 1070 9191 1104
rect 9191 1070 9225 1104
rect 9225 1070 9228 1104
rect 9176 1061 9228 1070
rect 9241 1104 9293 1113
rect 9306 1104 9358 1113
rect 9241 1070 9263 1104
rect 9263 1070 9293 1104
rect 9306 1070 9335 1104
rect 9335 1070 9358 1104
rect 9241 1061 9293 1070
rect 9306 1061 9358 1070
rect 9371 1061 9423 1113
rect 9436 1061 9488 1113
rect 9501 1104 9553 1113
rect 9566 1104 9618 1113
rect 9631 1104 9683 1113
rect 9696 1104 9748 1113
rect 9761 1104 9813 1113
rect 9826 1104 9878 1113
rect 9501 1070 9533 1104
rect 9533 1070 9553 1104
rect 9566 1070 9567 1104
rect 9567 1070 9605 1104
rect 9605 1070 9618 1104
rect 9631 1070 9639 1104
rect 9639 1070 9677 1104
rect 9677 1070 9683 1104
rect 9696 1070 9711 1104
rect 9711 1070 9748 1104
rect 9761 1070 9783 1104
rect 9783 1070 9813 1104
rect 9826 1070 9855 1104
rect 9855 1070 9878 1104
rect 9501 1061 9553 1070
rect 9566 1061 9618 1070
rect 9631 1061 9683 1070
rect 9696 1061 9748 1070
rect 9761 1061 9813 1070
rect 9826 1061 9878 1070
rect 9891 1104 9943 1113
rect 9891 1070 9893 1104
rect 9893 1070 9927 1104
rect 9927 1070 9943 1104
rect 9891 1061 9943 1070
rect 9956 1104 10008 1113
rect 9956 1070 9965 1104
rect 9965 1070 9999 1104
rect 9999 1070 10008 1104
rect 9956 1061 10008 1070
rect 10021 1104 10073 1113
rect 10021 1070 10037 1104
rect 10037 1070 10071 1104
rect 10071 1070 10073 1104
rect 10021 1061 10073 1070
rect 10086 1104 10138 1113
rect 10151 1104 10203 1113
rect 10216 1104 10268 1113
rect 10281 1104 10333 1113
rect 10346 1104 10398 1113
rect 10411 1104 10463 1113
rect 10476 1104 10528 1113
rect 10086 1070 10109 1104
rect 10109 1070 10138 1104
rect 10151 1070 10181 1104
rect 10181 1070 10203 1104
rect 10216 1070 10253 1104
rect 10253 1070 10268 1104
rect 10281 1070 10287 1104
rect 10287 1070 10325 1104
rect 10325 1070 10333 1104
rect 10346 1070 10359 1104
rect 10359 1070 10397 1104
rect 10397 1070 10398 1104
rect 10411 1070 10431 1104
rect 10431 1070 10463 1104
rect 10476 1070 10503 1104
rect 10503 1070 10528 1104
rect 10086 1061 10138 1070
rect 10151 1061 10203 1070
rect 10216 1061 10268 1070
rect 10281 1061 10333 1070
rect 10346 1061 10398 1070
rect 10411 1061 10463 1070
rect 10476 1061 10528 1070
rect 10541 1104 10593 1113
rect 10541 1070 10575 1104
rect 10575 1070 10593 1104
rect 10541 1061 10593 1070
rect 10606 1104 10658 1113
rect 10606 1070 10613 1104
rect 10613 1070 10647 1104
rect 10647 1070 10658 1104
rect 10606 1061 10658 1070
rect 10671 1104 10723 1113
rect 10671 1070 10685 1104
rect 10685 1070 10719 1104
rect 10719 1070 10723 1104
rect 10671 1061 10723 1070
rect 10736 1104 10788 1113
rect 10800 1104 10852 1113
rect 10864 1104 10916 1113
rect 10928 1104 10980 1113
rect 10992 1104 11044 1113
rect 11056 1104 11108 1113
rect 11120 1104 11172 1113
rect 10736 1070 10757 1104
rect 10757 1070 10788 1104
rect 10800 1070 10829 1104
rect 10829 1070 10852 1104
rect 10864 1070 10901 1104
rect 10901 1070 10916 1104
rect 10928 1070 10935 1104
rect 10935 1070 10973 1104
rect 10973 1070 10980 1104
rect 10992 1070 11007 1104
rect 11007 1070 11044 1104
rect 11056 1070 11079 1104
rect 11079 1070 11108 1104
rect 11120 1070 11151 1104
rect 11151 1070 11172 1104
rect 10736 1061 10788 1070
rect 10800 1061 10852 1070
rect 10864 1061 10916 1070
rect 10928 1061 10980 1070
rect 10992 1061 11044 1070
rect 11056 1061 11108 1070
rect 11120 1061 11172 1070
rect 11184 1104 11236 1113
rect 11184 1070 11189 1104
rect 11189 1070 11223 1104
rect 11223 1070 11236 1104
rect 11184 1061 11236 1070
rect 11248 1104 11300 1113
rect 11248 1070 11261 1104
rect 11261 1070 11295 1104
rect 11295 1070 11300 1104
rect 11248 1061 11300 1070
rect 11312 1104 11364 1113
rect 11376 1104 11428 1113
rect 11440 1104 11492 1113
rect 11504 1104 11556 1113
rect 11568 1104 11620 1113
rect 11632 1104 11684 1113
rect 11696 1104 11748 1113
rect 11312 1070 11333 1104
rect 11333 1070 11364 1104
rect 11376 1070 11405 1104
rect 11405 1070 11428 1104
rect 11440 1070 11477 1104
rect 11477 1070 11492 1104
rect 11504 1070 11511 1104
rect 11511 1070 11549 1104
rect 11549 1070 11556 1104
rect 11568 1070 11583 1104
rect 11583 1070 11620 1104
rect 11632 1070 11655 1104
rect 11655 1070 11684 1104
rect 11696 1070 11727 1104
rect 11727 1070 11748 1104
rect 11312 1061 11364 1070
rect 11376 1061 11428 1070
rect 11440 1061 11492 1070
rect 11504 1061 11556 1070
rect 11568 1061 11620 1070
rect 11632 1061 11684 1070
rect 11696 1061 11748 1070
rect 11760 1104 11812 1113
rect 11760 1070 11765 1104
rect 11765 1070 11799 1104
rect 11799 1070 11812 1104
rect 11760 1061 11812 1070
rect 11824 1104 11876 1113
rect 12022 1104 12074 1113
rect 12087 1104 12139 1113
rect 12152 1104 12204 1113
rect 12217 1104 12269 1113
rect 12282 1104 12334 1113
rect 12347 1104 12399 1113
rect 11824 1070 11837 1104
rect 11837 1070 11871 1104
rect 11871 1070 11876 1104
rect 12022 1070 12053 1104
rect 12053 1070 12074 1104
rect 12087 1070 12125 1104
rect 12125 1070 12139 1104
rect 12152 1070 12159 1104
rect 12159 1070 12197 1104
rect 12197 1070 12204 1104
rect 12217 1070 12231 1104
rect 12231 1070 12269 1104
rect 12282 1070 12303 1104
rect 12303 1070 12334 1104
rect 12347 1070 12375 1104
rect 12375 1070 12399 1104
rect 11824 1061 11876 1070
rect 12022 1061 12074 1070
rect 12087 1061 12139 1070
rect 12152 1061 12204 1070
rect 12217 1061 12269 1070
rect 12282 1061 12334 1070
rect 12347 1061 12399 1070
rect 12412 1104 12464 1113
rect 12412 1070 12413 1104
rect 12413 1070 12447 1104
rect 12447 1070 12464 1104
rect 12412 1061 12464 1070
rect 12477 1104 12529 1113
rect 12477 1070 12485 1104
rect 12485 1070 12519 1104
rect 12519 1070 12529 1104
rect 12477 1061 12529 1070
rect 12542 1061 12594 1113
rect 12607 1061 12659 1113
rect 12672 1104 12724 1113
rect 12672 1070 12683 1104
rect 12683 1070 12717 1104
rect 12717 1070 12724 1104
rect 12672 1061 12724 1070
rect 12737 1104 12789 1113
rect 12737 1070 12755 1104
rect 12755 1070 12789 1104
rect 12737 1061 12789 1070
rect 12801 1104 12853 1113
rect 12865 1104 12917 1113
rect 12929 1104 12981 1113
rect 12993 1104 13045 1113
rect 13057 1104 13109 1113
rect 13121 1104 13173 1113
rect 12801 1070 12827 1104
rect 12827 1070 12853 1104
rect 12865 1070 12899 1104
rect 12899 1070 12917 1104
rect 12929 1070 12933 1104
rect 12933 1070 12971 1104
rect 12971 1070 12981 1104
rect 12993 1070 13005 1104
rect 13005 1070 13043 1104
rect 13043 1070 13045 1104
rect 13057 1070 13077 1104
rect 13077 1070 13109 1104
rect 13121 1070 13149 1104
rect 13149 1070 13173 1104
rect 12801 1061 12853 1070
rect 12865 1061 12917 1070
rect 12929 1061 12981 1070
rect 12993 1061 13045 1070
rect 13057 1061 13109 1070
rect 13121 1061 13173 1070
rect 13185 1104 13237 1113
rect 13185 1070 13187 1104
rect 13187 1070 13221 1104
rect 13221 1070 13237 1104
rect 13185 1061 13237 1070
rect 13249 1104 13301 1113
rect 13249 1070 13259 1104
rect 13259 1070 13293 1104
rect 13293 1070 13301 1104
rect 13249 1061 13301 1070
rect 13313 1104 13365 1113
rect 13313 1070 13331 1104
rect 13331 1070 13365 1104
rect 13313 1061 13365 1070
rect 13377 1104 13429 1113
rect 13441 1104 13493 1113
rect 13505 1104 13557 1113
rect 13569 1104 13621 1113
rect 13633 1104 13685 1113
rect 13697 1104 13749 1113
rect 13377 1070 13403 1104
rect 13403 1070 13429 1104
rect 13441 1070 13475 1104
rect 13475 1070 13493 1104
rect 13505 1070 13509 1104
rect 13509 1070 13547 1104
rect 13547 1070 13557 1104
rect 13569 1070 13581 1104
rect 13581 1070 13619 1104
rect 13619 1070 13621 1104
rect 13633 1070 13653 1104
rect 13653 1070 13685 1104
rect 13697 1070 13725 1104
rect 13725 1070 13749 1104
rect 13377 1061 13429 1070
rect 13441 1061 13493 1070
rect 13505 1061 13557 1070
rect 13569 1061 13621 1070
rect 13633 1061 13685 1070
rect 13697 1061 13749 1070
rect 13761 1104 13813 1113
rect 13761 1070 13763 1104
rect 13763 1070 13797 1104
rect 13797 1070 13813 1104
rect 13761 1061 13813 1070
rect 13825 1104 13877 1113
rect 13825 1070 13835 1104
rect 13835 1070 13869 1104
rect 13869 1070 13877 1104
rect 13825 1061 13877 1070
rect 13889 1104 13941 1113
rect 13889 1070 13907 1104
rect 13907 1070 13941 1104
rect 13889 1061 13941 1070
rect 13953 1104 14005 1113
rect 14017 1104 14069 1113
rect 14081 1104 14133 1113
rect 14145 1104 14197 1113
rect 14209 1104 14261 1113
rect 14273 1104 14325 1113
rect 13953 1070 13979 1104
rect 13979 1070 14005 1104
rect 14017 1070 14051 1104
rect 14051 1070 14069 1104
rect 14081 1070 14085 1104
rect 14085 1070 14123 1104
rect 14123 1070 14133 1104
rect 14145 1070 14157 1104
rect 14157 1070 14195 1104
rect 14195 1070 14197 1104
rect 14209 1070 14229 1104
rect 14229 1070 14261 1104
rect 14273 1070 14301 1104
rect 14301 1070 14325 1104
rect 13953 1061 14005 1070
rect 14017 1061 14069 1070
rect 14081 1061 14133 1070
rect 14145 1061 14197 1070
rect 14209 1061 14261 1070
rect 14273 1061 14325 1070
rect 14337 1104 14389 1113
rect 14337 1070 14339 1104
rect 14339 1070 14373 1104
rect 14373 1070 14389 1104
rect 14337 1061 14389 1070
rect 14401 1104 14453 1113
rect 14401 1070 14411 1104
rect 14411 1070 14445 1104
rect 14445 1070 14453 1104
rect 14401 1061 14453 1070
rect 14465 1104 14517 1113
rect 14465 1070 14483 1104
rect 14483 1070 14517 1104
rect 14465 1061 14517 1070
rect 14529 1104 14581 1113
rect 14593 1104 14645 1113
rect 14657 1104 14709 1113
rect 14721 1104 14773 1113
rect 14785 1104 14837 1113
rect 14849 1104 14901 1113
rect 14529 1070 14555 1104
rect 14555 1070 14581 1104
rect 14593 1070 14627 1104
rect 14627 1070 14645 1104
rect 14657 1070 14661 1104
rect 14661 1070 14699 1104
rect 14699 1070 14709 1104
rect 14721 1070 14733 1104
rect 14733 1070 14771 1104
rect 14771 1070 14773 1104
rect 14785 1070 14805 1104
rect 14805 1070 14837 1104
rect 14849 1070 14877 1104
rect 14877 1070 14901 1104
rect 14529 1061 14581 1070
rect 14593 1061 14645 1070
rect 14657 1061 14709 1070
rect 14721 1061 14773 1070
rect 14785 1061 14837 1070
rect 14849 1061 14901 1070
rect 14913 1104 14965 1113
rect 14913 1070 14915 1104
rect 14915 1070 14949 1104
rect 14949 1070 14965 1104
rect 14913 1061 14965 1070
rect 14977 1104 15029 1113
rect 14977 1070 14987 1104
rect 14987 1070 15021 1104
rect 15021 1070 15029 1104
rect 14977 1061 15029 1070
rect 15041 1104 15093 1113
rect 15041 1070 15059 1104
rect 15059 1070 15093 1104
rect 15041 1061 15093 1070
rect 15105 1104 15157 1113
rect 15169 1104 15221 1113
rect 15233 1104 15285 1113
rect 15297 1104 15349 1113
rect 15361 1104 15413 1113
rect 15425 1104 15477 1113
rect 15105 1070 15131 1104
rect 15131 1070 15157 1104
rect 15169 1070 15203 1104
rect 15203 1070 15221 1104
rect 15233 1070 15237 1104
rect 15237 1070 15275 1104
rect 15275 1070 15285 1104
rect 15297 1070 15309 1104
rect 15309 1070 15347 1104
rect 15347 1070 15349 1104
rect 15361 1070 15381 1104
rect 15381 1070 15413 1104
rect 15425 1070 15453 1104
rect 15453 1070 15477 1104
rect 15105 1061 15157 1070
rect 15169 1061 15221 1070
rect 15233 1061 15285 1070
rect 15297 1061 15349 1070
rect 15361 1061 15413 1070
rect 15425 1061 15477 1070
rect 15489 1104 15541 1113
rect 15489 1070 15491 1104
rect 15491 1070 15525 1104
rect 15525 1070 15541 1104
rect 15489 1061 15541 1070
rect 15553 1104 15605 1113
rect 15553 1070 15563 1104
rect 15563 1070 15597 1104
rect 15597 1070 15605 1104
rect 15553 1061 15605 1070
rect 15617 1104 15669 1113
rect 15617 1070 15635 1104
rect 15635 1070 15669 1104
rect 15617 1061 15669 1070
rect 15681 1061 15733 1113
rect 15745 1061 15797 1113
rect 15809 1104 15861 1113
rect 15873 1104 15925 1113
rect 15937 1104 15989 1113
rect 16001 1104 16053 1113
rect 16065 1104 16117 1113
rect 16129 1104 16181 1113
rect 15809 1070 15833 1104
rect 15833 1070 15861 1104
rect 15873 1070 15905 1104
rect 15905 1070 15925 1104
rect 15937 1070 15939 1104
rect 15939 1070 15977 1104
rect 15977 1070 15989 1104
rect 16001 1070 16011 1104
rect 16011 1070 16049 1104
rect 16049 1070 16053 1104
rect 16065 1070 16083 1104
rect 16083 1070 16117 1104
rect 16129 1070 16155 1104
rect 16155 1070 16181 1104
rect 15809 1061 15861 1070
rect 15873 1061 15925 1070
rect 15937 1061 15989 1070
rect 16001 1061 16053 1070
rect 16065 1061 16117 1070
rect 16129 1061 16181 1070
rect 16193 1104 16245 1113
rect 16193 1070 16227 1104
rect 16227 1070 16245 1104
rect 16193 1061 16245 1070
rect 16257 1104 16309 1113
rect 16257 1070 16265 1104
rect 16265 1070 16299 1104
rect 16299 1070 16309 1104
rect 16257 1061 16309 1070
rect 16321 1104 16373 1113
rect 16321 1070 16337 1104
rect 16337 1070 16371 1104
rect 16371 1070 16373 1104
rect 16321 1061 16373 1070
rect 16385 1104 16437 1113
rect 16449 1104 16501 1113
rect 16513 1104 16565 1113
rect 16577 1104 16629 1113
rect 16641 1104 16693 1113
rect 16705 1104 16757 1113
rect 16385 1070 16409 1104
rect 16409 1070 16437 1104
rect 16449 1070 16481 1104
rect 16481 1070 16501 1104
rect 16513 1070 16515 1104
rect 16515 1070 16553 1104
rect 16553 1070 16565 1104
rect 16577 1070 16587 1104
rect 16587 1070 16625 1104
rect 16625 1070 16629 1104
rect 16641 1070 16659 1104
rect 16659 1070 16693 1104
rect 16705 1070 16731 1104
rect 16731 1070 16757 1104
rect 16385 1061 16437 1070
rect 16449 1061 16501 1070
rect 16513 1061 16565 1070
rect 16577 1061 16629 1070
rect 16641 1061 16693 1070
rect 16705 1061 16757 1070
rect 16769 1104 16821 1113
rect 16769 1070 16803 1104
rect 16803 1070 16821 1104
rect 16769 1061 16821 1070
rect 16833 1104 16885 1113
rect 16833 1070 16841 1104
rect 16841 1070 16875 1104
rect 16875 1070 16885 1104
rect 16833 1061 16885 1070
rect 16897 1104 16949 1113
rect 16897 1070 16913 1104
rect 16913 1070 16947 1104
rect 16947 1070 16949 1104
rect 16897 1061 16949 1070
rect 16961 1104 17013 1113
rect 17025 1104 17077 1113
rect 17089 1104 17141 1113
rect 17153 1104 17205 1113
rect 17217 1104 17269 1113
rect 17281 1104 17333 1113
rect 16961 1070 16985 1104
rect 16985 1070 17013 1104
rect 17025 1070 17057 1104
rect 17057 1070 17077 1104
rect 17089 1070 17091 1104
rect 17091 1070 17129 1104
rect 17129 1070 17141 1104
rect 17153 1070 17163 1104
rect 17163 1070 17201 1104
rect 17201 1070 17205 1104
rect 17217 1070 17235 1104
rect 17235 1070 17269 1104
rect 17281 1070 17307 1104
rect 17307 1070 17333 1104
rect 16961 1061 17013 1070
rect 17025 1061 17077 1070
rect 17089 1061 17141 1070
rect 17153 1061 17205 1070
rect 17217 1061 17269 1070
rect 17281 1061 17333 1070
rect 17345 1104 17397 1113
rect 17345 1070 17379 1104
rect 17379 1070 17397 1104
rect 17345 1061 17397 1070
rect 17409 1104 17461 1113
rect 17409 1070 17417 1104
rect 17417 1070 17451 1104
rect 17451 1070 17461 1104
rect 17409 1061 17461 1070
rect 17473 1104 17525 1113
rect 17473 1070 17489 1104
rect 17489 1070 17523 1104
rect 17523 1070 17525 1104
rect 17473 1061 17525 1070
rect 17537 1104 17589 1113
rect 17601 1104 17653 1113
rect 17665 1104 17717 1113
rect 17729 1104 17781 1113
rect 17793 1104 17845 1113
rect 17857 1104 17909 1113
rect 17537 1070 17561 1104
rect 17561 1070 17589 1104
rect 17601 1070 17633 1104
rect 17633 1070 17653 1104
rect 17665 1070 17667 1104
rect 17667 1070 17705 1104
rect 17705 1070 17717 1104
rect 17729 1070 17739 1104
rect 17739 1070 17777 1104
rect 17777 1070 17781 1104
rect 17793 1070 17811 1104
rect 17811 1070 17845 1104
rect 17857 1070 17883 1104
rect 17883 1070 17909 1104
rect 17537 1061 17589 1070
rect 17601 1061 17653 1070
rect 17665 1061 17717 1070
rect 17729 1061 17781 1070
rect 17793 1061 17845 1070
rect 17857 1061 17909 1070
rect 17921 1104 17973 1113
rect 17921 1070 17955 1104
rect 17955 1070 17973 1104
rect 17921 1061 17973 1070
rect 17985 1104 18037 1113
rect 17985 1070 17993 1104
rect 17993 1070 18027 1104
rect 18027 1070 18037 1104
rect 17985 1061 18037 1070
rect 18049 1104 18101 1113
rect 18049 1070 18065 1104
rect 18065 1070 18099 1104
rect 18099 1070 18101 1104
rect 18049 1061 18101 1070
rect 18113 1104 18165 1113
rect 18177 1104 18229 1113
rect 18241 1104 18293 1113
rect 18305 1104 18357 1113
rect 18369 1104 18421 1113
rect 18433 1104 18485 1113
rect 18113 1070 18137 1104
rect 18137 1070 18165 1104
rect 18177 1070 18209 1104
rect 18209 1070 18229 1104
rect 18241 1070 18243 1104
rect 18243 1070 18281 1104
rect 18281 1070 18293 1104
rect 18305 1070 18315 1104
rect 18315 1070 18353 1104
rect 18353 1070 18357 1104
rect 18369 1070 18387 1104
rect 18387 1070 18421 1104
rect 18433 1070 18459 1104
rect 18459 1070 18485 1104
rect 18113 1061 18165 1070
rect 18177 1061 18229 1070
rect 18241 1061 18293 1070
rect 18305 1061 18357 1070
rect 18369 1061 18421 1070
rect 18433 1061 18485 1070
rect 18497 1104 18549 1113
rect 18497 1070 18531 1104
rect 18531 1070 18549 1104
rect 18497 1061 18549 1070
rect 18561 1104 18613 1113
rect 18561 1070 18569 1104
rect 18569 1070 18603 1104
rect 18603 1070 18613 1104
rect 18561 1061 18613 1070
rect 18625 1104 18677 1113
rect 18625 1070 18641 1104
rect 18641 1070 18675 1104
rect 18675 1070 18677 1104
rect 18625 1061 18677 1070
rect 18689 1104 18741 1113
rect 18753 1104 18805 1113
rect 18817 1104 18869 1113
rect 18689 1070 18713 1104
rect 18713 1070 18741 1104
rect 18753 1070 18785 1104
rect 18785 1070 18805 1104
rect 18817 1070 18819 1104
rect 18819 1070 18869 1104
rect 18689 1061 18741 1070
rect 18753 1061 18805 1070
rect 18817 1061 18869 1070
rect 18881 1061 18933 1113
rect 18945 1104 18997 1113
rect 19009 1104 19061 1113
rect 19073 1104 19125 1113
rect 19137 1104 19189 1113
rect 19201 1104 19253 1113
rect 18945 1070 18983 1104
rect 18983 1070 18997 1104
rect 19009 1070 19017 1104
rect 19017 1070 19055 1104
rect 19055 1070 19061 1104
rect 19073 1070 19089 1104
rect 19089 1070 19125 1104
rect 19137 1070 19161 1104
rect 19161 1070 19189 1104
rect 19201 1070 19233 1104
rect 19233 1070 19253 1104
rect 18945 1061 18997 1070
rect 19009 1061 19061 1070
rect 19073 1061 19125 1070
rect 19137 1061 19189 1070
rect 19201 1061 19253 1070
rect 19265 1104 19317 1113
rect 19265 1070 19271 1104
rect 19271 1070 19305 1104
rect 19305 1070 19317 1104
rect 19265 1061 19317 1070
rect 19329 1104 19381 1113
rect 19329 1070 19343 1104
rect 19343 1070 19377 1104
rect 19377 1070 19381 1104
rect 19329 1061 19381 1070
rect 19393 1104 19445 1113
rect 19457 1104 19509 1113
rect 19521 1104 19573 1113
rect 19585 1104 19637 1113
rect 19649 1104 19701 1113
rect 19713 1104 19765 1113
rect 19777 1104 19829 1113
rect 19393 1070 19415 1104
rect 19415 1070 19445 1104
rect 19457 1070 19487 1104
rect 19487 1070 19509 1104
rect 19521 1070 19559 1104
rect 19559 1070 19573 1104
rect 19585 1070 19593 1104
rect 19593 1070 19631 1104
rect 19631 1070 19637 1104
rect 19649 1070 19665 1104
rect 19665 1070 19701 1104
rect 19713 1070 19737 1104
rect 19737 1070 19765 1104
rect 19777 1070 19809 1104
rect 19809 1070 19829 1104
rect 19393 1061 19445 1070
rect 19457 1061 19509 1070
rect 19521 1061 19573 1070
rect 19585 1061 19637 1070
rect 19649 1061 19701 1070
rect 19713 1061 19765 1070
rect 19777 1061 19829 1070
rect 19841 1104 19893 1113
rect 19841 1070 19847 1104
rect 19847 1070 19881 1104
rect 19881 1070 19893 1104
rect 19841 1061 19893 1070
rect 19905 1104 19957 1113
rect 19905 1070 19919 1104
rect 19919 1070 19953 1104
rect 19953 1070 19957 1104
rect 19905 1061 19957 1070
rect 19969 1104 20021 1113
rect 20033 1104 20085 1113
rect 20097 1104 20149 1113
rect 20161 1104 20213 1113
rect 20225 1104 20277 1113
rect 20289 1104 20341 1113
rect 20353 1104 20405 1113
rect 19969 1070 19991 1104
rect 19991 1070 20021 1104
rect 20033 1070 20063 1104
rect 20063 1070 20085 1104
rect 20097 1070 20135 1104
rect 20135 1070 20149 1104
rect 20161 1070 20169 1104
rect 20169 1070 20207 1104
rect 20207 1070 20213 1104
rect 20225 1070 20241 1104
rect 20241 1070 20277 1104
rect 20289 1070 20313 1104
rect 20313 1070 20341 1104
rect 20353 1070 20385 1104
rect 20385 1070 20405 1104
rect 19969 1061 20021 1070
rect 20033 1061 20085 1070
rect 20097 1061 20149 1070
rect 20161 1061 20213 1070
rect 20225 1061 20277 1070
rect 20289 1061 20341 1070
rect 20353 1061 20405 1070
rect 20417 1104 20469 1113
rect 20417 1070 20423 1104
rect 20423 1070 20457 1104
rect 20457 1070 20469 1104
rect 20417 1061 20469 1070
rect 20481 1104 20533 1113
rect 20481 1070 20495 1104
rect 20495 1070 20529 1104
rect 20529 1070 20533 1104
rect 20481 1061 20533 1070
rect 20545 1104 20597 1113
rect 20609 1104 20661 1113
rect 20673 1104 20725 1113
rect 20737 1104 20789 1113
rect 20801 1104 20853 1113
rect 20865 1104 20917 1113
rect 20929 1104 20981 1113
rect 20545 1070 20567 1104
rect 20567 1070 20597 1104
rect 20609 1070 20639 1104
rect 20639 1070 20661 1104
rect 20673 1070 20711 1104
rect 20711 1070 20725 1104
rect 20737 1070 20745 1104
rect 20745 1070 20783 1104
rect 20783 1070 20789 1104
rect 20801 1070 20817 1104
rect 20817 1070 20853 1104
rect 20865 1070 20889 1104
rect 20889 1070 20917 1104
rect 20929 1070 20961 1104
rect 20961 1070 20981 1104
rect 20545 1061 20597 1070
rect 20609 1061 20661 1070
rect 20673 1061 20725 1070
rect 20737 1061 20789 1070
rect 20801 1061 20853 1070
rect 20865 1061 20917 1070
rect 20929 1061 20981 1070
rect 20993 1104 21045 1113
rect 20993 1070 20999 1104
rect 20999 1070 21033 1104
rect 21033 1070 21045 1104
rect 20993 1061 21045 1070
rect 21057 1104 21109 1113
rect 21057 1070 21071 1104
rect 21071 1070 21105 1104
rect 21105 1070 21109 1104
rect 21057 1061 21109 1070
rect 21121 1104 21173 1113
rect 21185 1104 21237 1113
rect 21249 1104 21301 1113
rect 21313 1104 21365 1113
rect 21377 1104 21429 1113
rect 21441 1104 21493 1113
rect 21505 1104 21557 1113
rect 21121 1070 21143 1104
rect 21143 1070 21173 1104
rect 21185 1070 21215 1104
rect 21215 1070 21237 1104
rect 21249 1070 21287 1104
rect 21287 1070 21301 1104
rect 21313 1070 21321 1104
rect 21321 1070 21359 1104
rect 21359 1070 21365 1104
rect 21377 1070 21393 1104
rect 21393 1070 21429 1104
rect 21441 1070 21465 1104
rect 21465 1070 21493 1104
rect 21505 1070 21537 1104
rect 21537 1070 21557 1104
rect 21121 1061 21173 1070
rect 21185 1061 21237 1070
rect 21249 1061 21301 1070
rect 21313 1061 21365 1070
rect 21377 1061 21429 1070
rect 21441 1061 21493 1070
rect 21505 1061 21557 1070
rect 21569 1104 21621 1113
rect 21569 1070 21575 1104
rect 21575 1070 21609 1104
rect 21609 1070 21621 1104
rect 21569 1061 21621 1070
rect 21633 1104 21685 1113
rect 21633 1070 21647 1104
rect 21647 1070 21681 1104
rect 21681 1070 21685 1104
rect 21633 1061 21685 1070
rect 21697 1104 21749 1113
rect 21761 1104 21813 1113
rect 21825 1104 21877 1113
rect 21889 1104 21941 1113
rect 21697 1070 21719 1104
rect 21719 1070 21749 1104
rect 21761 1070 21791 1104
rect 21791 1070 21813 1104
rect 21825 1070 21863 1104
rect 21863 1070 21877 1104
rect 21889 1070 21897 1104
rect 21897 1070 21935 1104
rect 21935 1070 21941 1104
rect 21697 1061 21749 1070
rect 21761 1061 21813 1070
rect 21825 1061 21877 1070
rect 21889 1061 21941 1070
rect 22236 1107 22248 1140
rect 22248 1107 22282 1140
rect 22282 1107 22288 1140
rect 22439 1170 22491 1179
rect 22439 1136 22472 1170
rect 22472 1136 22491 1170
rect 22439 1127 22491 1136
rect 22507 1170 22559 1179
rect 22507 1136 22510 1170
rect 22510 1136 22544 1170
rect 22544 1136 22559 1170
rect 22507 1127 22559 1136
rect 22575 1170 22627 1179
rect 22575 1136 22582 1170
rect 22582 1136 22616 1170
rect 22616 1136 22627 1170
rect 22575 1127 22627 1136
rect 22643 1170 22695 1179
rect 22643 1136 22654 1170
rect 22654 1136 22688 1170
rect 22688 1136 22695 1170
rect 22643 1127 22695 1136
rect 22711 1170 22763 1179
rect 22711 1136 22726 1170
rect 22726 1136 22760 1170
rect 22760 1136 22763 1170
rect 22711 1127 22763 1136
rect 22779 1170 22831 1179
rect 22847 1170 22899 1179
rect 22915 1170 22967 1179
rect 22982 1170 23034 1179
rect 23049 1170 23101 1179
rect 23116 1170 23168 1179
rect 23183 1170 23235 1179
rect 23250 1170 23302 1179
rect 22779 1136 22798 1170
rect 22798 1136 22831 1170
rect 22847 1136 22870 1170
rect 22870 1136 22899 1170
rect 22915 1136 22942 1170
rect 22942 1136 22967 1170
rect 22982 1136 23014 1170
rect 23014 1136 23034 1170
rect 23049 1136 23086 1170
rect 23086 1136 23101 1170
rect 23116 1136 23120 1170
rect 23120 1136 23158 1170
rect 23158 1136 23168 1170
rect 23183 1136 23192 1170
rect 23192 1136 23230 1170
rect 23230 1136 23235 1170
rect 23250 1136 23264 1170
rect 23264 1136 23302 1170
rect 22779 1127 22831 1136
rect 22847 1127 22899 1136
rect 22915 1127 22967 1136
rect 22982 1127 23034 1136
rect 23049 1127 23101 1136
rect 23116 1127 23168 1136
rect 23183 1127 23235 1136
rect 23250 1127 23302 1136
rect 22236 1064 22288 1095
rect 22236 1043 22248 1064
rect 22248 1043 22282 1064
rect 22282 1043 22288 1064
rect 22236 1030 22248 1031
rect 22248 1030 22282 1031
rect 22282 1030 22288 1031
rect 22236 988 22288 1030
rect 22236 979 22248 988
rect 22248 979 22282 988
rect 22282 979 22288 988
rect 23407 1014 23459 1022
rect 23478 1014 23530 1022
rect 23549 1014 23601 1022
rect 23620 1014 23672 1022
rect 23691 1014 23743 1022
rect 23762 1014 23814 1022
rect 23833 1014 23885 1022
rect 23904 1014 23956 1022
rect 23975 1014 24027 1022
rect 24046 1014 24098 1022
rect 23407 980 23408 1014
rect 23408 980 23446 1014
rect 23446 980 23459 1014
rect 23478 980 23480 1014
rect 23480 980 23518 1014
rect 23518 980 23530 1014
rect 23549 980 23552 1014
rect 23552 980 23590 1014
rect 23590 980 23601 1014
rect 23620 980 23624 1014
rect 23624 980 23662 1014
rect 23662 980 23672 1014
rect 23691 980 23696 1014
rect 23696 980 23734 1014
rect 23734 980 23743 1014
rect 23762 980 23768 1014
rect 23768 980 23806 1014
rect 23806 980 23814 1014
rect 23833 980 23840 1014
rect 23840 980 23878 1014
rect 23878 980 23885 1014
rect 23904 980 23912 1014
rect 23912 980 23950 1014
rect 23950 980 23956 1014
rect 23975 980 23984 1014
rect 23984 980 24022 1014
rect 24022 980 24027 1014
rect 24046 980 24056 1014
rect 24056 980 24094 1014
rect 24094 980 24098 1014
rect 23407 970 23459 980
rect 23478 970 23530 980
rect 23549 970 23601 980
rect 23620 970 23672 980
rect 23691 970 23743 980
rect 23762 970 23814 980
rect 23833 970 23885 980
rect 23904 970 23956 980
rect 23975 970 24027 980
rect 24046 970 24098 980
rect 7616 948 7668 957
rect 7681 948 7733 957
rect 7616 914 7641 948
rect 7641 914 7668 948
rect 7681 914 7713 948
rect 7713 914 7733 948
rect 7616 905 7668 914
rect 7681 905 7733 914
rect 7746 948 7798 957
rect 7746 914 7751 948
rect 7751 914 7785 948
rect 7785 914 7798 948
rect 7746 905 7798 914
rect 7811 948 7863 957
rect 7811 914 7823 948
rect 7823 914 7857 948
rect 7857 914 7863 948
rect 7811 905 7863 914
rect 7876 948 7928 957
rect 7941 948 7993 957
rect 8006 948 8058 957
rect 8071 948 8123 957
rect 8136 948 8188 957
rect 8201 948 8253 957
rect 8266 948 8318 957
rect 8331 948 8383 957
rect 7876 914 7895 948
rect 7895 914 7928 948
rect 7941 914 7967 948
rect 7967 914 7993 948
rect 8006 914 8039 948
rect 8039 914 8058 948
rect 8071 914 8073 948
rect 8073 914 8111 948
rect 8111 914 8123 948
rect 8136 914 8145 948
rect 8145 914 8183 948
rect 8183 914 8188 948
rect 8201 914 8217 948
rect 8217 914 8253 948
rect 8266 914 8289 948
rect 8289 914 8318 948
rect 8331 914 8361 948
rect 8361 914 8383 948
rect 7876 905 7928 914
rect 7941 905 7993 914
rect 8006 905 8058 914
rect 8071 905 8123 914
rect 8136 905 8188 914
rect 8201 905 8253 914
rect 8266 905 8318 914
rect 8331 905 8383 914
rect 8396 948 8448 957
rect 8396 914 8399 948
rect 8399 914 8433 948
rect 8433 914 8448 948
rect 8396 905 8448 914
rect 8461 948 8513 957
rect 8461 914 8471 948
rect 8471 914 8505 948
rect 8505 914 8513 948
rect 8461 905 8513 914
rect 8526 948 8578 957
rect 8526 914 8543 948
rect 8543 914 8577 948
rect 8577 914 8578 948
rect 8526 905 8578 914
rect 8591 948 8643 957
rect 8656 948 8708 957
rect 8721 948 8773 957
rect 8786 948 8838 957
rect 8851 948 8903 957
rect 8916 948 8968 957
rect 8981 948 9033 957
rect 8591 914 8615 948
rect 8615 914 8643 948
rect 8656 914 8687 948
rect 8687 914 8708 948
rect 8721 914 8759 948
rect 8759 914 8773 948
rect 8786 914 8793 948
rect 8793 914 8831 948
rect 8831 914 8838 948
rect 8851 914 8865 948
rect 8865 914 8903 948
rect 8916 914 8937 948
rect 8937 914 8968 948
rect 8981 914 9009 948
rect 9009 914 9033 948
rect 8591 905 8643 914
rect 8656 905 8708 914
rect 8721 905 8773 914
rect 8786 905 8838 914
rect 8851 905 8903 914
rect 8916 905 8968 914
rect 8981 905 9033 914
rect 9046 948 9098 957
rect 9046 914 9047 948
rect 9047 914 9081 948
rect 9081 914 9098 948
rect 9046 905 9098 914
rect 9111 948 9163 957
rect 9111 914 9119 948
rect 9119 914 9153 948
rect 9153 914 9163 948
rect 9111 905 9163 914
rect 9176 948 9228 957
rect 9176 914 9191 948
rect 9191 914 9225 948
rect 9225 914 9228 948
rect 9176 905 9228 914
rect 9241 948 9293 957
rect 9306 948 9358 957
rect 9241 914 9263 948
rect 9263 914 9293 948
rect 9306 914 9335 948
rect 9335 914 9358 948
rect 9241 905 9293 914
rect 9306 905 9358 914
rect 9371 905 9423 957
rect 9436 905 9488 957
rect 9501 948 9553 957
rect 9566 948 9618 957
rect 9631 948 9683 957
rect 9696 948 9748 957
rect 9761 948 9813 957
rect 9826 948 9878 957
rect 9501 914 9533 948
rect 9533 914 9553 948
rect 9566 914 9567 948
rect 9567 914 9605 948
rect 9605 914 9618 948
rect 9631 914 9639 948
rect 9639 914 9677 948
rect 9677 914 9683 948
rect 9696 914 9711 948
rect 9711 914 9748 948
rect 9761 914 9783 948
rect 9783 914 9813 948
rect 9826 914 9855 948
rect 9855 914 9878 948
rect 9501 905 9553 914
rect 9566 905 9618 914
rect 9631 905 9683 914
rect 9696 905 9748 914
rect 9761 905 9813 914
rect 9826 905 9878 914
rect 9891 948 9943 957
rect 9891 914 9893 948
rect 9893 914 9927 948
rect 9927 914 9943 948
rect 9891 905 9943 914
rect 9956 948 10008 957
rect 9956 914 9965 948
rect 9965 914 9999 948
rect 9999 914 10008 948
rect 9956 905 10008 914
rect 10021 948 10073 957
rect 10021 914 10037 948
rect 10037 914 10071 948
rect 10071 914 10073 948
rect 10021 905 10073 914
rect 10086 948 10138 957
rect 10151 948 10203 957
rect 10216 948 10268 957
rect 10281 948 10333 957
rect 10346 948 10398 957
rect 10411 948 10463 957
rect 10476 948 10528 957
rect 10086 914 10109 948
rect 10109 914 10138 948
rect 10151 914 10181 948
rect 10181 914 10203 948
rect 10216 914 10253 948
rect 10253 914 10268 948
rect 10281 914 10287 948
rect 10287 914 10325 948
rect 10325 914 10333 948
rect 10346 914 10359 948
rect 10359 914 10397 948
rect 10397 914 10398 948
rect 10411 914 10431 948
rect 10431 914 10463 948
rect 10476 914 10503 948
rect 10503 914 10528 948
rect 10086 905 10138 914
rect 10151 905 10203 914
rect 10216 905 10268 914
rect 10281 905 10333 914
rect 10346 905 10398 914
rect 10411 905 10463 914
rect 10476 905 10528 914
rect 10541 948 10593 957
rect 10541 914 10575 948
rect 10575 914 10593 948
rect 10541 905 10593 914
rect 10606 948 10658 957
rect 10606 914 10613 948
rect 10613 914 10647 948
rect 10647 914 10658 948
rect 10606 905 10658 914
rect 10671 948 10723 957
rect 10671 914 10685 948
rect 10685 914 10719 948
rect 10719 914 10723 948
rect 10671 905 10723 914
rect 10736 948 10788 957
rect 10800 948 10852 957
rect 10864 948 10916 957
rect 10928 948 10980 957
rect 10992 948 11044 957
rect 11056 948 11108 957
rect 11120 948 11172 957
rect 10736 914 10757 948
rect 10757 914 10788 948
rect 10800 914 10829 948
rect 10829 914 10852 948
rect 10864 914 10901 948
rect 10901 914 10916 948
rect 10928 914 10935 948
rect 10935 914 10973 948
rect 10973 914 10980 948
rect 10992 914 11007 948
rect 11007 914 11044 948
rect 11056 914 11079 948
rect 11079 914 11108 948
rect 11120 914 11151 948
rect 11151 914 11172 948
rect 10736 905 10788 914
rect 10800 905 10852 914
rect 10864 905 10916 914
rect 10928 905 10980 914
rect 10992 905 11044 914
rect 11056 905 11108 914
rect 11120 905 11172 914
rect 11184 948 11236 957
rect 11184 914 11189 948
rect 11189 914 11223 948
rect 11223 914 11236 948
rect 11184 905 11236 914
rect 11248 948 11300 957
rect 11248 914 11261 948
rect 11261 914 11295 948
rect 11295 914 11300 948
rect 11248 905 11300 914
rect 11312 948 11364 957
rect 11376 948 11428 957
rect 11440 948 11492 957
rect 11504 948 11556 957
rect 11568 948 11620 957
rect 11632 948 11684 957
rect 11696 948 11748 957
rect 11312 914 11333 948
rect 11333 914 11364 948
rect 11376 914 11405 948
rect 11405 914 11428 948
rect 11440 914 11477 948
rect 11477 914 11492 948
rect 11504 914 11511 948
rect 11511 914 11549 948
rect 11549 914 11556 948
rect 11568 914 11583 948
rect 11583 914 11620 948
rect 11632 914 11655 948
rect 11655 914 11684 948
rect 11696 914 11727 948
rect 11727 914 11748 948
rect 11312 905 11364 914
rect 11376 905 11428 914
rect 11440 905 11492 914
rect 11504 905 11556 914
rect 11568 905 11620 914
rect 11632 905 11684 914
rect 11696 905 11748 914
rect 11760 948 11812 957
rect 11760 914 11765 948
rect 11765 914 11799 948
rect 11799 914 11812 948
rect 11760 905 11812 914
rect 11824 948 11876 957
rect 12022 948 12074 957
rect 12087 948 12139 957
rect 12152 948 12204 957
rect 12217 948 12269 957
rect 12282 948 12334 957
rect 12347 948 12399 957
rect 11824 914 11837 948
rect 11837 914 11871 948
rect 11871 914 11876 948
rect 12022 914 12053 948
rect 12053 914 12074 948
rect 12087 914 12125 948
rect 12125 914 12139 948
rect 12152 914 12159 948
rect 12159 914 12197 948
rect 12197 914 12204 948
rect 12217 914 12231 948
rect 12231 914 12269 948
rect 12282 914 12303 948
rect 12303 914 12334 948
rect 12347 914 12375 948
rect 12375 914 12399 948
rect 11824 905 11876 914
rect 12022 905 12074 914
rect 12087 905 12139 914
rect 12152 905 12204 914
rect 12217 905 12269 914
rect 12282 905 12334 914
rect 12347 905 12399 914
rect 12412 948 12464 957
rect 12412 914 12413 948
rect 12413 914 12447 948
rect 12447 914 12464 948
rect 12412 905 12464 914
rect 12477 948 12529 957
rect 12477 914 12485 948
rect 12485 914 12519 948
rect 12519 914 12529 948
rect 12477 905 12529 914
rect 12542 905 12594 957
rect 12607 905 12659 957
rect 12672 948 12724 957
rect 12672 914 12683 948
rect 12683 914 12717 948
rect 12717 914 12724 948
rect 12672 905 12724 914
rect 12737 948 12789 957
rect 12737 914 12755 948
rect 12755 914 12789 948
rect 12737 905 12789 914
rect 12802 948 12854 957
rect 12867 948 12919 957
rect 12932 948 12984 957
rect 12997 948 13049 957
rect 13062 948 13114 957
rect 13127 948 13179 957
rect 13192 948 13244 957
rect 12802 914 12827 948
rect 12827 914 12854 948
rect 12867 914 12899 948
rect 12899 914 12919 948
rect 12932 914 12933 948
rect 12933 914 12971 948
rect 12971 914 12984 948
rect 12997 914 13005 948
rect 13005 914 13043 948
rect 13043 914 13049 948
rect 13062 914 13077 948
rect 13077 914 13114 948
rect 13127 914 13149 948
rect 13149 914 13179 948
rect 13192 914 13221 948
rect 13221 914 13244 948
rect 12802 905 12854 914
rect 12867 905 12919 914
rect 12932 905 12984 914
rect 12997 905 13049 914
rect 13062 905 13114 914
rect 13127 905 13179 914
rect 13192 905 13244 914
rect 13257 948 13309 957
rect 13257 914 13259 948
rect 13259 914 13293 948
rect 13293 914 13309 948
rect 13257 905 13309 914
rect 13322 948 13374 957
rect 13322 914 13331 948
rect 13331 914 13365 948
rect 13365 914 13374 948
rect 13322 905 13374 914
rect 13387 948 13439 957
rect 13387 914 13403 948
rect 13403 914 13437 948
rect 13437 914 13439 948
rect 13387 905 13439 914
rect 13452 948 13504 957
rect 13517 948 13569 957
rect 13582 948 13634 957
rect 13647 948 13699 957
rect 13712 948 13764 957
rect 13777 948 13829 957
rect 13842 948 13894 957
rect 13452 914 13475 948
rect 13475 914 13504 948
rect 13517 914 13547 948
rect 13547 914 13569 948
rect 13582 914 13619 948
rect 13619 914 13634 948
rect 13647 914 13653 948
rect 13653 914 13691 948
rect 13691 914 13699 948
rect 13712 914 13725 948
rect 13725 914 13763 948
rect 13763 914 13764 948
rect 13777 914 13797 948
rect 13797 914 13829 948
rect 13842 914 13869 948
rect 13869 914 13894 948
rect 13452 905 13504 914
rect 13517 905 13569 914
rect 13582 905 13634 914
rect 13647 905 13699 914
rect 13712 905 13764 914
rect 13777 905 13829 914
rect 13842 905 13894 914
rect 13907 948 13959 957
rect 13907 914 13941 948
rect 13941 914 13959 948
rect 13907 905 13959 914
rect 13972 948 14024 957
rect 13972 914 13979 948
rect 13979 914 14013 948
rect 14013 914 14024 948
rect 13972 905 14024 914
rect 14037 948 14089 957
rect 14037 914 14051 948
rect 14051 914 14085 948
rect 14085 914 14089 948
rect 14037 905 14089 914
rect 14102 948 14154 957
rect 14167 948 14219 957
rect 14232 948 14284 957
rect 14297 948 14349 957
rect 14362 948 14414 957
rect 14427 948 14479 957
rect 14492 948 14544 957
rect 14557 948 14609 957
rect 14102 914 14123 948
rect 14123 914 14154 948
rect 14167 914 14195 948
rect 14195 914 14219 948
rect 14232 914 14267 948
rect 14267 914 14284 948
rect 14297 914 14301 948
rect 14301 914 14339 948
rect 14339 914 14349 948
rect 14362 914 14373 948
rect 14373 914 14411 948
rect 14411 914 14414 948
rect 14427 914 14445 948
rect 14445 914 14479 948
rect 14492 914 14517 948
rect 14517 914 14544 948
rect 14557 914 14589 948
rect 14589 914 14609 948
rect 14102 905 14154 914
rect 14167 905 14219 914
rect 14232 905 14284 914
rect 14297 905 14349 914
rect 14362 905 14414 914
rect 14427 905 14479 914
rect 14492 905 14544 914
rect 14557 905 14609 914
rect 14622 948 14674 957
rect 14622 914 14627 948
rect 14627 914 14661 948
rect 14661 914 14674 948
rect 14622 905 14674 914
rect 14686 948 14738 957
rect 14686 914 14699 948
rect 14699 914 14733 948
rect 14733 914 14738 948
rect 14686 905 14738 914
rect 14750 948 14802 957
rect 14814 948 14866 957
rect 14878 948 14930 957
rect 14942 948 14994 957
rect 15006 948 15058 957
rect 15070 948 15122 957
rect 15134 948 15186 957
rect 14750 914 14771 948
rect 14771 914 14802 948
rect 14814 914 14843 948
rect 14843 914 14866 948
rect 14878 914 14915 948
rect 14915 914 14930 948
rect 14942 914 14949 948
rect 14949 914 14987 948
rect 14987 914 14994 948
rect 15006 914 15021 948
rect 15021 914 15058 948
rect 15070 914 15093 948
rect 15093 914 15122 948
rect 15134 914 15165 948
rect 15165 914 15186 948
rect 14750 905 14802 914
rect 14814 905 14866 914
rect 14878 905 14930 914
rect 14942 905 14994 914
rect 15006 905 15058 914
rect 15070 905 15122 914
rect 15134 905 15186 914
rect 15198 948 15250 957
rect 15198 914 15203 948
rect 15203 914 15237 948
rect 15237 914 15250 948
rect 15198 905 15250 914
rect 15262 948 15314 957
rect 15262 914 15275 948
rect 15275 914 15309 948
rect 15309 914 15314 948
rect 15262 905 15314 914
rect 15326 948 15378 957
rect 15390 948 15442 957
rect 15454 948 15506 957
rect 15518 948 15570 957
rect 15582 948 15634 957
rect 15646 948 15698 957
rect 15326 914 15347 948
rect 15347 914 15378 948
rect 15390 914 15419 948
rect 15419 914 15442 948
rect 15454 914 15491 948
rect 15491 914 15506 948
rect 15518 914 15525 948
rect 15525 914 15563 948
rect 15563 914 15570 948
rect 15582 914 15597 948
rect 15597 914 15634 948
rect 15646 914 15669 948
rect 15669 914 15698 948
rect 15326 905 15378 914
rect 15390 905 15442 914
rect 15454 905 15506 914
rect 15518 905 15570 914
rect 15582 905 15634 914
rect 15646 905 15698 914
rect 15710 905 15762 957
rect 15774 905 15826 957
rect 15838 948 15890 957
rect 15838 914 15867 948
rect 15867 914 15890 948
rect 15838 905 15890 914
rect 15902 948 15954 957
rect 15902 914 15905 948
rect 15905 914 15939 948
rect 15939 914 15954 948
rect 15902 905 15954 914
rect 15966 948 16018 957
rect 15966 914 15977 948
rect 15977 914 16011 948
rect 16011 914 16018 948
rect 15966 905 16018 914
rect 16030 948 16082 957
rect 16094 948 16146 957
rect 16158 948 16210 957
rect 16222 948 16274 957
rect 16286 948 16338 957
rect 16350 948 16402 957
rect 16414 948 16466 957
rect 16030 914 16049 948
rect 16049 914 16082 948
rect 16094 914 16121 948
rect 16121 914 16146 948
rect 16158 914 16193 948
rect 16193 914 16210 948
rect 16222 914 16227 948
rect 16227 914 16265 948
rect 16265 914 16274 948
rect 16286 914 16299 948
rect 16299 914 16337 948
rect 16337 914 16338 948
rect 16350 914 16371 948
rect 16371 914 16402 948
rect 16414 914 16443 948
rect 16443 914 16466 948
rect 16030 905 16082 914
rect 16094 905 16146 914
rect 16158 905 16210 914
rect 16222 905 16274 914
rect 16286 905 16338 914
rect 16350 905 16402 914
rect 16414 905 16466 914
rect 16478 948 16530 957
rect 16478 914 16481 948
rect 16481 914 16515 948
rect 16515 914 16530 948
rect 16478 905 16530 914
rect 16542 948 16594 957
rect 16542 914 16553 948
rect 16553 914 16587 948
rect 16587 914 16594 948
rect 16542 905 16594 914
rect 16606 948 16658 957
rect 16670 948 16722 957
rect 16734 948 16786 957
rect 16798 948 16850 957
rect 16862 948 16914 957
rect 16926 948 16978 957
rect 16990 948 17042 957
rect 16606 914 16625 948
rect 16625 914 16658 948
rect 16670 914 16697 948
rect 16697 914 16722 948
rect 16734 914 16769 948
rect 16769 914 16786 948
rect 16798 914 16803 948
rect 16803 914 16841 948
rect 16841 914 16850 948
rect 16862 914 16875 948
rect 16875 914 16913 948
rect 16913 914 16914 948
rect 16926 914 16947 948
rect 16947 914 16978 948
rect 16990 914 17019 948
rect 17019 914 17042 948
rect 16606 905 16658 914
rect 16670 905 16722 914
rect 16734 905 16786 914
rect 16798 905 16850 914
rect 16862 905 16914 914
rect 16926 905 16978 914
rect 16990 905 17042 914
rect 17054 948 17106 957
rect 17054 914 17057 948
rect 17057 914 17091 948
rect 17091 914 17106 948
rect 17054 905 17106 914
rect 17118 948 17170 957
rect 17118 914 17129 948
rect 17129 914 17163 948
rect 17163 914 17170 948
rect 17118 905 17170 914
rect 17182 948 17234 957
rect 17246 948 17298 957
rect 17310 948 17362 957
rect 17374 948 17426 957
rect 17438 948 17490 957
rect 17502 948 17554 957
rect 17566 948 17618 957
rect 17182 914 17201 948
rect 17201 914 17234 948
rect 17246 914 17273 948
rect 17273 914 17298 948
rect 17310 914 17345 948
rect 17345 914 17362 948
rect 17374 914 17379 948
rect 17379 914 17417 948
rect 17417 914 17426 948
rect 17438 914 17451 948
rect 17451 914 17489 948
rect 17489 914 17490 948
rect 17502 914 17523 948
rect 17523 914 17554 948
rect 17566 914 17595 948
rect 17595 914 17618 948
rect 17182 905 17234 914
rect 17246 905 17298 914
rect 17310 905 17362 914
rect 17374 905 17426 914
rect 17438 905 17490 914
rect 17502 905 17554 914
rect 17566 905 17618 914
rect 17630 948 17682 957
rect 17630 914 17633 948
rect 17633 914 17667 948
rect 17667 914 17682 948
rect 17630 905 17682 914
rect 17694 948 17746 957
rect 17694 914 17705 948
rect 17705 914 17739 948
rect 17739 914 17746 948
rect 17694 905 17746 914
rect 17758 948 17810 957
rect 17822 948 17874 957
rect 17886 948 17938 957
rect 17950 948 18002 957
rect 18014 948 18066 957
rect 18078 948 18130 957
rect 18142 948 18194 957
rect 17758 914 17777 948
rect 17777 914 17810 948
rect 17822 914 17849 948
rect 17849 914 17874 948
rect 17886 914 17921 948
rect 17921 914 17938 948
rect 17950 914 17955 948
rect 17955 914 17993 948
rect 17993 914 18002 948
rect 18014 914 18027 948
rect 18027 914 18065 948
rect 18065 914 18066 948
rect 18078 914 18099 948
rect 18099 914 18130 948
rect 18142 914 18171 948
rect 18171 914 18194 948
rect 17758 905 17810 914
rect 17822 905 17874 914
rect 17886 905 17938 914
rect 17950 905 18002 914
rect 18014 905 18066 914
rect 18078 905 18130 914
rect 18142 905 18194 914
rect 18206 948 18258 957
rect 18206 914 18209 948
rect 18209 914 18243 948
rect 18243 914 18258 948
rect 18206 905 18258 914
rect 18270 948 18322 957
rect 18270 914 18281 948
rect 18281 914 18315 948
rect 18315 914 18322 948
rect 18270 905 18322 914
rect 18334 948 18386 957
rect 18398 948 18450 957
rect 18462 948 18514 957
rect 18526 948 18578 957
rect 18590 948 18642 957
rect 18654 948 18706 957
rect 18718 948 18770 957
rect 18334 914 18353 948
rect 18353 914 18386 948
rect 18398 914 18425 948
rect 18425 914 18450 948
rect 18462 914 18497 948
rect 18497 914 18514 948
rect 18526 914 18531 948
rect 18531 914 18569 948
rect 18569 914 18578 948
rect 18590 914 18603 948
rect 18603 914 18641 948
rect 18641 914 18642 948
rect 18654 914 18675 948
rect 18675 914 18706 948
rect 18718 914 18747 948
rect 18747 914 18770 948
rect 18334 905 18386 914
rect 18398 905 18450 914
rect 18462 905 18514 914
rect 18526 905 18578 914
rect 18590 905 18642 914
rect 18654 905 18706 914
rect 18718 905 18770 914
rect 18782 948 18834 957
rect 18782 914 18785 948
rect 18785 914 18819 948
rect 18819 914 18834 948
rect 18782 905 18834 914
rect 18846 905 18898 957
rect 18910 905 18962 957
rect 18974 948 19026 957
rect 18974 914 18983 948
rect 18983 914 19017 948
rect 19017 914 19026 948
rect 18974 905 19026 914
rect 19038 948 19090 957
rect 19038 914 19055 948
rect 19055 914 19089 948
rect 19089 914 19090 948
rect 19038 905 19090 914
rect 19102 948 19154 957
rect 19166 948 19218 957
rect 19230 948 19282 957
rect 19294 948 19346 957
rect 19358 948 19410 957
rect 19422 948 19474 957
rect 19102 914 19127 948
rect 19127 914 19154 948
rect 19166 914 19199 948
rect 19199 914 19218 948
rect 19230 914 19233 948
rect 19233 914 19271 948
rect 19271 914 19282 948
rect 19294 914 19305 948
rect 19305 914 19343 948
rect 19343 914 19346 948
rect 19358 914 19377 948
rect 19377 914 19410 948
rect 19422 914 19449 948
rect 19449 914 19474 948
rect 19102 905 19154 914
rect 19166 905 19218 914
rect 19230 905 19282 914
rect 19294 905 19346 914
rect 19358 905 19410 914
rect 19422 905 19474 914
rect 19486 948 19538 957
rect 19486 914 19487 948
rect 19487 914 19521 948
rect 19521 914 19538 948
rect 19486 905 19538 914
rect 19550 948 19602 957
rect 19550 914 19559 948
rect 19559 914 19593 948
rect 19593 914 19602 948
rect 19550 905 19602 914
rect 19614 948 19666 957
rect 19614 914 19631 948
rect 19631 914 19665 948
rect 19665 914 19666 948
rect 19614 905 19666 914
rect 19678 948 19730 957
rect 19742 948 19794 957
rect 19806 948 19858 957
rect 19870 948 19922 957
rect 19934 948 19986 957
rect 19998 948 20050 957
rect 19678 914 19703 948
rect 19703 914 19730 948
rect 19742 914 19775 948
rect 19775 914 19794 948
rect 19806 914 19809 948
rect 19809 914 19847 948
rect 19847 914 19858 948
rect 19870 914 19881 948
rect 19881 914 19919 948
rect 19919 914 19922 948
rect 19934 914 19953 948
rect 19953 914 19986 948
rect 19998 914 20025 948
rect 20025 914 20050 948
rect 19678 905 19730 914
rect 19742 905 19794 914
rect 19806 905 19858 914
rect 19870 905 19922 914
rect 19934 905 19986 914
rect 19998 905 20050 914
rect 20062 948 20114 957
rect 20062 914 20063 948
rect 20063 914 20097 948
rect 20097 914 20114 948
rect 20062 905 20114 914
rect 20126 948 20178 957
rect 20126 914 20135 948
rect 20135 914 20169 948
rect 20169 914 20178 948
rect 20126 905 20178 914
rect 20190 948 20242 957
rect 20190 914 20207 948
rect 20207 914 20241 948
rect 20241 914 20242 948
rect 20190 905 20242 914
rect 20254 948 20306 957
rect 20318 948 20370 957
rect 20382 948 20434 957
rect 20446 948 20498 957
rect 20510 948 20562 957
rect 20574 948 20626 957
rect 20254 914 20279 948
rect 20279 914 20306 948
rect 20318 914 20351 948
rect 20351 914 20370 948
rect 20382 914 20385 948
rect 20385 914 20423 948
rect 20423 914 20434 948
rect 20446 914 20457 948
rect 20457 914 20495 948
rect 20495 914 20498 948
rect 20510 914 20529 948
rect 20529 914 20562 948
rect 20574 914 20601 948
rect 20601 914 20626 948
rect 20254 905 20306 914
rect 20318 905 20370 914
rect 20382 905 20434 914
rect 20446 905 20498 914
rect 20510 905 20562 914
rect 20574 905 20626 914
rect 20638 948 20690 957
rect 20638 914 20639 948
rect 20639 914 20673 948
rect 20673 914 20690 948
rect 20638 905 20690 914
rect 20702 948 20754 957
rect 20702 914 20711 948
rect 20711 914 20745 948
rect 20745 914 20754 948
rect 20702 905 20754 914
rect 20766 948 20818 957
rect 20766 914 20783 948
rect 20783 914 20817 948
rect 20817 914 20818 948
rect 20766 905 20818 914
rect 20830 948 20882 957
rect 20894 948 20946 957
rect 20958 948 21010 957
rect 21022 948 21074 957
rect 21086 948 21138 957
rect 21150 948 21202 957
rect 20830 914 20855 948
rect 20855 914 20882 948
rect 20894 914 20927 948
rect 20927 914 20946 948
rect 20958 914 20961 948
rect 20961 914 20999 948
rect 20999 914 21010 948
rect 21022 914 21033 948
rect 21033 914 21071 948
rect 21071 914 21074 948
rect 21086 914 21105 948
rect 21105 914 21138 948
rect 21150 914 21177 948
rect 21177 914 21202 948
rect 20830 905 20882 914
rect 20894 905 20946 914
rect 20958 905 21010 914
rect 21022 905 21074 914
rect 21086 905 21138 914
rect 21150 905 21202 914
rect 21214 948 21266 957
rect 21214 914 21215 948
rect 21215 914 21249 948
rect 21249 914 21266 948
rect 21214 905 21266 914
rect 21278 948 21330 957
rect 21278 914 21287 948
rect 21287 914 21321 948
rect 21321 914 21330 948
rect 21278 905 21330 914
rect 21342 948 21394 957
rect 21342 914 21359 948
rect 21359 914 21393 948
rect 21393 914 21394 948
rect 21342 905 21394 914
rect 21406 948 21458 957
rect 21470 948 21522 957
rect 21534 948 21586 957
rect 21598 948 21650 957
rect 21662 948 21714 957
rect 21726 948 21778 957
rect 21406 914 21431 948
rect 21431 914 21458 948
rect 21470 914 21503 948
rect 21503 914 21522 948
rect 21534 914 21537 948
rect 21537 914 21575 948
rect 21575 914 21586 948
rect 21598 914 21609 948
rect 21609 914 21647 948
rect 21647 914 21650 948
rect 21662 914 21681 948
rect 21681 914 21714 948
rect 21726 914 21753 948
rect 21753 914 21778 948
rect 21406 905 21458 914
rect 21470 905 21522 914
rect 21534 905 21586 914
rect 21598 905 21650 914
rect 21662 905 21714 914
rect 21726 905 21778 914
rect 21790 948 21842 957
rect 21790 914 21791 948
rect 21791 914 21825 948
rect 21825 914 21842 948
rect 21790 905 21842 914
rect 21854 948 21906 957
rect 21854 914 21863 948
rect 21863 914 21897 948
rect 21897 914 21906 948
rect 21854 905 21906 914
rect 21918 948 21970 957
rect 21918 914 21935 948
rect 21935 914 21969 948
rect 21969 914 21970 948
rect 21918 905 21970 914
rect 22236 954 22248 967
rect 22248 954 22282 967
rect 22282 954 22288 967
rect 22236 915 22288 954
rect 22236 878 22248 902
rect 22248 878 22282 902
rect 22282 878 22288 902
rect 22236 850 22288 878
rect 22236 836 22288 837
rect 1545 818 1597 827
rect 1610 818 1662 827
rect 1675 818 1727 827
rect 1740 818 1792 827
rect 1545 784 1557 818
rect 1557 784 1595 818
rect 1595 784 1597 818
rect 1610 784 1629 818
rect 1629 784 1662 818
rect 1675 784 1701 818
rect 1701 784 1727 818
rect 1740 784 1773 818
rect 1773 784 1792 818
rect 1545 775 1597 784
rect 1610 775 1662 784
rect 1675 775 1727 784
rect 1740 775 1792 784
rect 1805 818 1857 827
rect 1805 784 1811 818
rect 1811 784 1845 818
rect 1845 784 1857 818
rect 1805 775 1857 784
rect 1870 818 1922 827
rect 1870 784 1883 818
rect 1883 784 1917 818
rect 1917 784 1922 818
rect 1870 775 1922 784
rect 1935 818 1987 827
rect 2000 818 2052 827
rect 2065 818 2117 827
rect 2130 818 2182 827
rect 2195 818 2247 827
rect 2260 818 2312 827
rect 2325 818 2377 827
rect 2390 818 2442 827
rect 1935 784 1955 818
rect 1955 784 1987 818
rect 2000 784 2027 818
rect 2027 784 2052 818
rect 2065 784 2099 818
rect 2099 784 2117 818
rect 2130 784 2133 818
rect 2133 784 2171 818
rect 2171 784 2182 818
rect 2195 784 2205 818
rect 2205 784 2243 818
rect 2243 784 2247 818
rect 2260 784 2277 818
rect 2277 784 2312 818
rect 2325 784 2349 818
rect 2349 784 2377 818
rect 2390 784 2421 818
rect 2421 784 2442 818
rect 1935 775 1987 784
rect 2000 775 2052 784
rect 2065 775 2117 784
rect 2130 775 2182 784
rect 2195 775 2247 784
rect 2260 775 2312 784
rect 2325 775 2377 784
rect 2390 775 2442 784
rect 2455 818 2507 827
rect 2455 784 2459 818
rect 2459 784 2493 818
rect 2493 784 2507 818
rect 2455 775 2507 784
rect 2520 818 2572 827
rect 2520 784 2531 818
rect 2531 784 2565 818
rect 2565 784 2572 818
rect 2520 775 2572 784
rect 2585 818 2637 827
rect 2585 784 2603 818
rect 2603 784 2637 818
rect 2585 775 2637 784
rect 2650 818 2702 827
rect 2715 818 2767 827
rect 2780 818 2832 827
rect 2845 818 2897 827
rect 2910 818 2962 827
rect 2975 818 3027 827
rect 3040 818 3092 827
rect 2650 784 2675 818
rect 2675 784 2702 818
rect 2715 784 2747 818
rect 2747 784 2767 818
rect 2780 784 2781 818
rect 2781 784 2819 818
rect 2819 784 2832 818
rect 2845 784 2853 818
rect 2853 784 2891 818
rect 2891 784 2897 818
rect 2910 784 2925 818
rect 2925 784 2962 818
rect 2975 784 2997 818
rect 2997 784 3027 818
rect 3040 784 3069 818
rect 3069 784 3092 818
rect 2650 775 2702 784
rect 2715 775 2767 784
rect 2780 775 2832 784
rect 2845 775 2897 784
rect 2910 775 2962 784
rect 2975 775 3027 784
rect 3040 775 3092 784
rect 3105 775 3157 827
rect 3170 775 3222 827
rect 3235 818 3287 827
rect 3235 784 3267 818
rect 3267 784 3287 818
rect 3235 775 3287 784
rect 3300 818 3352 827
rect 3300 784 3305 818
rect 3305 784 3339 818
rect 3339 784 3352 818
rect 3300 775 3352 784
rect 3365 818 3417 827
rect 3365 784 3377 818
rect 3377 784 3411 818
rect 3411 784 3417 818
rect 3365 775 3417 784
rect 3430 818 3482 827
rect 3495 818 3547 827
rect 3560 818 3612 827
rect 3625 818 3677 827
rect 3690 818 3742 827
rect 3755 818 3807 827
rect 3820 818 3872 827
rect 3885 818 3937 827
rect 3430 784 3449 818
rect 3449 784 3482 818
rect 3495 784 3521 818
rect 3521 784 3547 818
rect 3560 784 3593 818
rect 3593 784 3612 818
rect 3625 784 3627 818
rect 3627 784 3665 818
rect 3665 784 3677 818
rect 3690 784 3699 818
rect 3699 784 3737 818
rect 3737 784 3742 818
rect 3755 784 3771 818
rect 3771 784 3807 818
rect 3820 784 3843 818
rect 3843 784 3872 818
rect 3885 784 3915 818
rect 3915 784 3937 818
rect 3430 775 3482 784
rect 3495 775 3547 784
rect 3560 775 3612 784
rect 3625 775 3677 784
rect 3690 775 3742 784
rect 3755 775 3807 784
rect 3820 775 3872 784
rect 3885 775 3937 784
rect 3950 818 4002 827
rect 3950 784 3953 818
rect 3953 784 3987 818
rect 3987 784 4002 818
rect 3950 775 4002 784
rect 4015 818 4067 827
rect 4015 784 4025 818
rect 4025 784 4059 818
rect 4059 784 4067 818
rect 4015 775 4067 784
rect 4080 818 4132 827
rect 4080 784 4097 818
rect 4097 784 4131 818
rect 4131 784 4132 818
rect 4080 775 4132 784
rect 4144 818 4196 827
rect 4208 818 4260 827
rect 4272 818 4324 827
rect 4336 818 4388 827
rect 4400 818 4452 827
rect 4464 818 4516 827
rect 4144 784 4169 818
rect 4169 784 4196 818
rect 4208 784 4241 818
rect 4241 784 4260 818
rect 4272 784 4275 818
rect 4275 784 4313 818
rect 4313 784 4324 818
rect 4336 784 4347 818
rect 4347 784 4385 818
rect 4385 784 4388 818
rect 4400 784 4419 818
rect 4419 784 4452 818
rect 4464 784 4491 818
rect 4491 784 4516 818
rect 4144 775 4196 784
rect 4208 775 4260 784
rect 4272 775 4324 784
rect 4336 775 4388 784
rect 4400 775 4452 784
rect 4464 775 4516 784
rect 4528 818 4580 827
rect 4528 784 4529 818
rect 4529 784 4563 818
rect 4563 784 4580 818
rect 4528 775 4580 784
rect 4592 818 4644 827
rect 4592 784 4601 818
rect 4601 784 4635 818
rect 4635 784 4644 818
rect 4592 775 4644 784
rect 4656 818 4708 827
rect 4656 784 4673 818
rect 4673 784 4707 818
rect 4707 784 4708 818
rect 4656 775 4708 784
rect 4720 818 4772 827
rect 4784 818 4836 827
rect 4848 818 4900 827
rect 4912 818 4964 827
rect 4976 818 5028 827
rect 5040 818 5092 827
rect 4720 784 4745 818
rect 4745 784 4772 818
rect 4784 784 4817 818
rect 4817 784 4836 818
rect 4848 784 4851 818
rect 4851 784 4889 818
rect 4889 784 4900 818
rect 4912 784 4923 818
rect 4923 784 4961 818
rect 4961 784 4964 818
rect 4976 784 4995 818
rect 4995 784 5028 818
rect 5040 784 5067 818
rect 5067 784 5092 818
rect 4720 775 4772 784
rect 4784 775 4836 784
rect 4848 775 4900 784
rect 4912 775 4964 784
rect 4976 775 5028 784
rect 5040 775 5092 784
rect 5104 818 5156 827
rect 5104 784 5105 818
rect 5105 784 5139 818
rect 5139 784 5156 818
rect 5104 775 5156 784
rect 5168 818 5220 827
rect 5168 784 5177 818
rect 5177 784 5211 818
rect 5211 784 5220 818
rect 5168 775 5220 784
rect 5232 818 5284 827
rect 5232 784 5249 818
rect 5249 784 5283 818
rect 5283 784 5284 818
rect 5232 775 5284 784
rect 5296 818 5348 827
rect 5360 818 5412 827
rect 5424 818 5476 827
rect 5488 818 5540 827
rect 5552 818 5604 827
rect 5616 818 5668 827
rect 5296 784 5321 818
rect 5321 784 5348 818
rect 5360 784 5393 818
rect 5393 784 5412 818
rect 5424 784 5427 818
rect 5427 784 5465 818
rect 5465 784 5476 818
rect 5488 784 5499 818
rect 5499 784 5537 818
rect 5537 784 5540 818
rect 5552 784 5571 818
rect 5571 784 5604 818
rect 5616 784 5643 818
rect 5643 784 5668 818
rect 5296 775 5348 784
rect 5360 775 5412 784
rect 5424 775 5476 784
rect 5488 775 5540 784
rect 5552 775 5604 784
rect 5616 775 5668 784
rect 5680 818 5732 827
rect 5680 784 5681 818
rect 5681 784 5715 818
rect 5715 784 5732 818
rect 5680 775 5732 784
rect 5744 818 5796 827
rect 5744 784 5753 818
rect 5753 784 5787 818
rect 5787 784 5796 818
rect 5744 775 5796 784
rect 5808 818 5860 827
rect 5808 784 5825 818
rect 5825 784 5859 818
rect 5859 784 5860 818
rect 5808 775 5860 784
rect 5872 818 5924 827
rect 5936 818 5988 827
rect 6000 818 6052 827
rect 6064 818 6116 827
rect 5872 784 5897 818
rect 5897 784 5924 818
rect 5936 784 5969 818
rect 5969 784 5988 818
rect 6000 784 6003 818
rect 6003 784 6041 818
rect 6041 784 6052 818
rect 6064 784 6075 818
rect 6075 784 6113 818
rect 6113 784 6116 818
rect 5872 775 5924 784
rect 5936 775 5988 784
rect 6000 775 6052 784
rect 6064 775 6116 784
rect 22236 802 22248 836
rect 22248 802 22282 836
rect 22282 802 22288 836
rect 22439 858 22491 867
rect 22439 824 22472 858
rect 22472 824 22491 858
rect 22439 815 22491 824
rect 22507 858 22559 867
rect 22507 824 22510 858
rect 22510 824 22544 858
rect 22544 824 22559 858
rect 22507 815 22559 824
rect 22575 858 22627 867
rect 22575 824 22582 858
rect 22582 824 22616 858
rect 22616 824 22627 858
rect 22575 815 22627 824
rect 22643 858 22695 867
rect 22643 824 22654 858
rect 22654 824 22688 858
rect 22688 824 22695 858
rect 22643 815 22695 824
rect 22711 858 22763 867
rect 22711 824 22726 858
rect 22726 824 22760 858
rect 22760 824 22763 858
rect 22711 815 22763 824
rect 22779 858 22831 867
rect 22847 858 22899 867
rect 22915 858 22967 867
rect 22982 858 23034 867
rect 23049 858 23101 867
rect 23116 858 23168 867
rect 23183 858 23235 867
rect 23250 858 23302 867
rect 22779 824 22798 858
rect 22798 824 22831 858
rect 22847 824 22870 858
rect 22870 824 22899 858
rect 22915 824 22942 858
rect 22942 824 22967 858
rect 22982 824 23014 858
rect 23014 824 23034 858
rect 23049 824 23086 858
rect 23086 824 23101 858
rect 23116 824 23120 858
rect 23120 824 23158 858
rect 23158 824 23168 858
rect 23183 824 23192 858
rect 23192 824 23230 858
rect 23230 824 23235 858
rect 23250 824 23264 858
rect 23264 824 23302 858
rect 22779 815 22831 824
rect 22847 815 22899 824
rect 22915 815 22967 824
rect 22982 815 23034 824
rect 23049 815 23101 824
rect 23116 815 23168 824
rect 23183 815 23235 824
rect 23250 815 23302 824
rect 7616 792 7668 801
rect 7681 792 7733 801
rect 7616 758 7641 792
rect 7641 758 7668 792
rect 7681 758 7713 792
rect 7713 758 7733 792
rect 7616 749 7668 758
rect 7681 749 7733 758
rect 7746 792 7798 801
rect 7746 758 7751 792
rect 7751 758 7785 792
rect 7785 758 7798 792
rect 7746 749 7798 758
rect 7811 792 7863 801
rect 7811 758 7823 792
rect 7823 758 7857 792
rect 7857 758 7863 792
rect 7811 749 7863 758
rect 7876 792 7928 801
rect 7941 792 7993 801
rect 8006 792 8058 801
rect 8071 792 8123 801
rect 8136 792 8188 801
rect 8201 792 8253 801
rect 8266 792 8318 801
rect 8331 792 8383 801
rect 7876 758 7895 792
rect 7895 758 7928 792
rect 7941 758 7967 792
rect 7967 758 7993 792
rect 8006 758 8039 792
rect 8039 758 8058 792
rect 8071 758 8073 792
rect 8073 758 8111 792
rect 8111 758 8123 792
rect 8136 758 8145 792
rect 8145 758 8183 792
rect 8183 758 8188 792
rect 8201 758 8217 792
rect 8217 758 8253 792
rect 8266 758 8289 792
rect 8289 758 8318 792
rect 8331 758 8361 792
rect 8361 758 8383 792
rect 7876 749 7928 758
rect 7941 749 7993 758
rect 8006 749 8058 758
rect 8071 749 8123 758
rect 8136 749 8188 758
rect 8201 749 8253 758
rect 8266 749 8318 758
rect 8331 749 8383 758
rect 8396 792 8448 801
rect 8396 758 8399 792
rect 8399 758 8433 792
rect 8433 758 8448 792
rect 8396 749 8448 758
rect 8461 792 8513 801
rect 8461 758 8471 792
rect 8471 758 8505 792
rect 8505 758 8513 792
rect 8461 749 8513 758
rect 8526 792 8578 801
rect 8526 758 8543 792
rect 8543 758 8577 792
rect 8577 758 8578 792
rect 8526 749 8578 758
rect 8591 792 8643 801
rect 8656 792 8708 801
rect 8721 792 8773 801
rect 8786 792 8838 801
rect 8851 792 8903 801
rect 8916 792 8968 801
rect 8981 792 9033 801
rect 8591 758 8615 792
rect 8615 758 8643 792
rect 8656 758 8687 792
rect 8687 758 8708 792
rect 8721 758 8759 792
rect 8759 758 8773 792
rect 8786 758 8793 792
rect 8793 758 8831 792
rect 8831 758 8838 792
rect 8851 758 8865 792
rect 8865 758 8903 792
rect 8916 758 8937 792
rect 8937 758 8968 792
rect 8981 758 9009 792
rect 9009 758 9033 792
rect 8591 749 8643 758
rect 8656 749 8708 758
rect 8721 749 8773 758
rect 8786 749 8838 758
rect 8851 749 8903 758
rect 8916 749 8968 758
rect 8981 749 9033 758
rect 9046 792 9098 801
rect 9046 758 9047 792
rect 9047 758 9081 792
rect 9081 758 9098 792
rect 9046 749 9098 758
rect 9111 792 9163 801
rect 9111 758 9119 792
rect 9119 758 9153 792
rect 9153 758 9163 792
rect 9111 749 9163 758
rect 9176 792 9228 801
rect 9176 758 9191 792
rect 9191 758 9225 792
rect 9225 758 9228 792
rect 9176 749 9228 758
rect 9241 792 9293 801
rect 9306 792 9358 801
rect 9241 758 9263 792
rect 9263 758 9293 792
rect 9306 758 9335 792
rect 9335 758 9358 792
rect 9241 749 9293 758
rect 9306 749 9358 758
rect 9371 749 9423 801
rect 9436 749 9488 801
rect 9501 792 9553 801
rect 9566 792 9618 801
rect 9631 792 9683 801
rect 9696 792 9748 801
rect 9761 792 9813 801
rect 9826 792 9878 801
rect 9501 758 9533 792
rect 9533 758 9553 792
rect 9566 758 9567 792
rect 9567 758 9605 792
rect 9605 758 9618 792
rect 9631 758 9639 792
rect 9639 758 9677 792
rect 9677 758 9683 792
rect 9696 758 9711 792
rect 9711 758 9748 792
rect 9761 758 9783 792
rect 9783 758 9813 792
rect 9826 758 9855 792
rect 9855 758 9878 792
rect 9501 749 9553 758
rect 9566 749 9618 758
rect 9631 749 9683 758
rect 9696 749 9748 758
rect 9761 749 9813 758
rect 9826 749 9878 758
rect 9891 792 9943 801
rect 9891 758 9893 792
rect 9893 758 9927 792
rect 9927 758 9943 792
rect 9891 749 9943 758
rect 9956 792 10008 801
rect 9956 758 9965 792
rect 9965 758 9999 792
rect 9999 758 10008 792
rect 9956 749 10008 758
rect 10021 792 10073 801
rect 10021 758 10037 792
rect 10037 758 10071 792
rect 10071 758 10073 792
rect 10021 749 10073 758
rect 10086 792 10138 801
rect 10151 792 10203 801
rect 10216 792 10268 801
rect 10281 792 10333 801
rect 10346 792 10398 801
rect 10411 792 10463 801
rect 10476 792 10528 801
rect 10086 758 10109 792
rect 10109 758 10138 792
rect 10151 758 10181 792
rect 10181 758 10203 792
rect 10216 758 10253 792
rect 10253 758 10268 792
rect 10281 758 10287 792
rect 10287 758 10325 792
rect 10325 758 10333 792
rect 10346 758 10359 792
rect 10359 758 10397 792
rect 10397 758 10398 792
rect 10411 758 10431 792
rect 10431 758 10463 792
rect 10476 758 10503 792
rect 10503 758 10528 792
rect 10086 749 10138 758
rect 10151 749 10203 758
rect 10216 749 10268 758
rect 10281 749 10333 758
rect 10346 749 10398 758
rect 10411 749 10463 758
rect 10476 749 10528 758
rect 10541 792 10593 801
rect 10541 758 10575 792
rect 10575 758 10593 792
rect 10541 749 10593 758
rect 10606 792 10658 801
rect 10606 758 10613 792
rect 10613 758 10647 792
rect 10647 758 10658 792
rect 10606 749 10658 758
rect 10671 792 10723 801
rect 10671 758 10685 792
rect 10685 758 10719 792
rect 10719 758 10723 792
rect 10671 749 10723 758
rect 10736 792 10788 801
rect 10800 792 10852 801
rect 10864 792 10916 801
rect 10928 792 10980 801
rect 10992 792 11044 801
rect 11056 792 11108 801
rect 11120 792 11172 801
rect 10736 758 10757 792
rect 10757 758 10788 792
rect 10800 758 10829 792
rect 10829 758 10852 792
rect 10864 758 10901 792
rect 10901 758 10916 792
rect 10928 758 10935 792
rect 10935 758 10973 792
rect 10973 758 10980 792
rect 10992 758 11007 792
rect 11007 758 11044 792
rect 11056 758 11079 792
rect 11079 758 11108 792
rect 11120 758 11151 792
rect 11151 758 11172 792
rect 10736 749 10788 758
rect 10800 749 10852 758
rect 10864 749 10916 758
rect 10928 749 10980 758
rect 10992 749 11044 758
rect 11056 749 11108 758
rect 11120 749 11172 758
rect 11184 792 11236 801
rect 11184 758 11189 792
rect 11189 758 11223 792
rect 11223 758 11236 792
rect 11184 749 11236 758
rect 11248 792 11300 801
rect 11248 758 11261 792
rect 11261 758 11295 792
rect 11295 758 11300 792
rect 11248 749 11300 758
rect 11312 792 11364 801
rect 11376 792 11428 801
rect 11440 792 11492 801
rect 11504 792 11556 801
rect 11568 792 11620 801
rect 11632 792 11684 801
rect 11696 792 11748 801
rect 11312 758 11333 792
rect 11333 758 11364 792
rect 11376 758 11405 792
rect 11405 758 11428 792
rect 11440 758 11477 792
rect 11477 758 11492 792
rect 11504 758 11511 792
rect 11511 758 11549 792
rect 11549 758 11556 792
rect 11568 758 11583 792
rect 11583 758 11620 792
rect 11632 758 11655 792
rect 11655 758 11684 792
rect 11696 758 11727 792
rect 11727 758 11748 792
rect 11312 749 11364 758
rect 11376 749 11428 758
rect 11440 749 11492 758
rect 11504 749 11556 758
rect 11568 749 11620 758
rect 11632 749 11684 758
rect 11696 749 11748 758
rect 11760 792 11812 801
rect 11760 758 11765 792
rect 11765 758 11799 792
rect 11799 758 11812 792
rect 11760 749 11812 758
rect 11824 792 11876 801
rect 12022 792 12074 801
rect 12087 792 12139 801
rect 12152 792 12204 801
rect 12217 792 12269 801
rect 12282 792 12334 801
rect 12347 792 12399 801
rect 11824 758 11837 792
rect 11837 758 11871 792
rect 11871 758 11876 792
rect 12022 758 12053 792
rect 12053 758 12074 792
rect 12087 758 12125 792
rect 12125 758 12139 792
rect 12152 758 12159 792
rect 12159 758 12197 792
rect 12197 758 12204 792
rect 12217 758 12231 792
rect 12231 758 12269 792
rect 12282 758 12303 792
rect 12303 758 12334 792
rect 12347 758 12375 792
rect 12375 758 12399 792
rect 11824 749 11876 758
rect 12022 749 12074 758
rect 12087 749 12139 758
rect 12152 749 12204 758
rect 12217 749 12269 758
rect 12282 749 12334 758
rect 12347 749 12399 758
rect 12412 792 12464 801
rect 12412 758 12413 792
rect 12413 758 12447 792
rect 12447 758 12464 792
rect 12412 749 12464 758
rect 12477 792 12529 801
rect 12477 758 12485 792
rect 12485 758 12519 792
rect 12519 758 12529 792
rect 12477 749 12529 758
rect 12542 749 12594 801
rect 12607 749 12659 801
rect 12672 792 12724 801
rect 12672 758 12683 792
rect 12683 758 12717 792
rect 12717 758 12724 792
rect 12672 749 12724 758
rect 12737 792 12789 801
rect 12737 758 12755 792
rect 12755 758 12789 792
rect 12737 749 12789 758
rect 12802 792 12854 801
rect 12867 792 12919 801
rect 12932 792 12984 801
rect 12997 792 13049 801
rect 13062 792 13114 801
rect 13127 792 13179 801
rect 13192 792 13244 801
rect 12802 758 12827 792
rect 12827 758 12854 792
rect 12867 758 12899 792
rect 12899 758 12919 792
rect 12932 758 12933 792
rect 12933 758 12971 792
rect 12971 758 12984 792
rect 12997 758 13005 792
rect 13005 758 13043 792
rect 13043 758 13049 792
rect 13062 758 13077 792
rect 13077 758 13114 792
rect 13127 758 13149 792
rect 13149 758 13179 792
rect 13192 758 13221 792
rect 13221 758 13244 792
rect 12802 749 12854 758
rect 12867 749 12919 758
rect 12932 749 12984 758
rect 12997 749 13049 758
rect 13062 749 13114 758
rect 13127 749 13179 758
rect 13192 749 13244 758
rect 13257 792 13309 801
rect 13257 758 13259 792
rect 13259 758 13293 792
rect 13293 758 13309 792
rect 13257 749 13309 758
rect 13322 792 13374 801
rect 13322 758 13331 792
rect 13331 758 13365 792
rect 13365 758 13374 792
rect 13322 749 13374 758
rect 13387 792 13439 801
rect 13387 758 13403 792
rect 13403 758 13437 792
rect 13437 758 13439 792
rect 13387 749 13439 758
rect 13452 792 13504 801
rect 13517 792 13569 801
rect 13582 792 13634 801
rect 13647 792 13699 801
rect 13712 792 13764 801
rect 13777 792 13829 801
rect 13842 792 13894 801
rect 13452 758 13475 792
rect 13475 758 13504 792
rect 13517 758 13547 792
rect 13547 758 13569 792
rect 13582 758 13619 792
rect 13619 758 13634 792
rect 13647 758 13653 792
rect 13653 758 13691 792
rect 13691 758 13699 792
rect 13712 758 13725 792
rect 13725 758 13763 792
rect 13763 758 13764 792
rect 13777 758 13797 792
rect 13797 758 13829 792
rect 13842 758 13869 792
rect 13869 758 13894 792
rect 13452 749 13504 758
rect 13517 749 13569 758
rect 13582 749 13634 758
rect 13647 749 13699 758
rect 13712 749 13764 758
rect 13777 749 13829 758
rect 13842 749 13894 758
rect 13907 792 13959 801
rect 13907 758 13941 792
rect 13941 758 13959 792
rect 13907 749 13959 758
rect 13972 792 14024 801
rect 13972 758 13979 792
rect 13979 758 14013 792
rect 14013 758 14024 792
rect 13972 749 14024 758
rect 14037 792 14089 801
rect 14037 758 14051 792
rect 14051 758 14085 792
rect 14085 758 14089 792
rect 14037 749 14089 758
rect 14101 792 14153 801
rect 14165 792 14217 801
rect 14229 792 14281 801
rect 14293 792 14345 801
rect 14357 792 14409 801
rect 14421 792 14473 801
rect 14485 792 14537 801
rect 14101 758 14123 792
rect 14123 758 14153 792
rect 14165 758 14195 792
rect 14195 758 14217 792
rect 14229 758 14267 792
rect 14267 758 14281 792
rect 14293 758 14301 792
rect 14301 758 14339 792
rect 14339 758 14345 792
rect 14357 758 14373 792
rect 14373 758 14409 792
rect 14421 758 14445 792
rect 14445 758 14473 792
rect 14485 758 14517 792
rect 14517 758 14537 792
rect 14101 749 14153 758
rect 14165 749 14217 758
rect 14229 749 14281 758
rect 14293 749 14345 758
rect 14357 749 14409 758
rect 14421 749 14473 758
rect 14485 749 14537 758
rect 14549 792 14601 801
rect 14549 758 14555 792
rect 14555 758 14589 792
rect 14589 758 14601 792
rect 14549 749 14601 758
rect 14613 792 14665 801
rect 14613 758 14627 792
rect 14627 758 14661 792
rect 14661 758 14665 792
rect 14613 749 14665 758
rect 14677 792 14729 801
rect 14741 792 14793 801
rect 14805 792 14857 801
rect 14869 792 14921 801
rect 14933 792 14985 801
rect 14997 792 15049 801
rect 15061 792 15113 801
rect 14677 758 14699 792
rect 14699 758 14729 792
rect 14741 758 14771 792
rect 14771 758 14793 792
rect 14805 758 14843 792
rect 14843 758 14857 792
rect 14869 758 14877 792
rect 14877 758 14915 792
rect 14915 758 14921 792
rect 14933 758 14949 792
rect 14949 758 14985 792
rect 14997 758 15021 792
rect 15021 758 15049 792
rect 15061 758 15093 792
rect 15093 758 15113 792
rect 14677 749 14729 758
rect 14741 749 14793 758
rect 14805 749 14857 758
rect 14869 749 14921 758
rect 14933 749 14985 758
rect 14997 749 15049 758
rect 15061 749 15113 758
rect 15125 792 15177 801
rect 15125 758 15131 792
rect 15131 758 15165 792
rect 15165 758 15177 792
rect 15125 749 15177 758
rect 15189 792 15241 801
rect 15189 758 15203 792
rect 15203 758 15237 792
rect 15237 758 15241 792
rect 15189 749 15241 758
rect 15253 792 15305 801
rect 15317 792 15369 801
rect 15381 792 15433 801
rect 15445 792 15497 801
rect 15509 792 15561 801
rect 15573 792 15625 801
rect 15637 792 15689 801
rect 15253 758 15275 792
rect 15275 758 15305 792
rect 15317 758 15347 792
rect 15347 758 15369 792
rect 15381 758 15419 792
rect 15419 758 15433 792
rect 15445 758 15453 792
rect 15453 758 15491 792
rect 15491 758 15497 792
rect 15509 758 15525 792
rect 15525 758 15561 792
rect 15573 758 15597 792
rect 15597 758 15625 792
rect 15637 758 15669 792
rect 15669 758 15689 792
rect 15253 749 15305 758
rect 15317 749 15369 758
rect 15381 749 15433 758
rect 15445 749 15497 758
rect 15509 749 15561 758
rect 15573 749 15625 758
rect 15637 749 15689 758
rect 15701 749 15753 801
rect 15765 749 15817 801
rect 15829 792 15881 801
rect 15829 758 15833 792
rect 15833 758 15867 792
rect 15867 758 15881 792
rect 15829 749 15881 758
rect 15893 792 15945 801
rect 15893 758 15905 792
rect 15905 758 15939 792
rect 15939 758 15945 792
rect 15893 749 15945 758
rect 15957 792 16009 801
rect 16021 792 16073 801
rect 16085 792 16137 801
rect 16149 792 16201 801
rect 16213 792 16265 801
rect 16277 792 16329 801
rect 16341 792 16393 801
rect 15957 758 15977 792
rect 15977 758 16009 792
rect 16021 758 16049 792
rect 16049 758 16073 792
rect 16085 758 16121 792
rect 16121 758 16137 792
rect 16149 758 16155 792
rect 16155 758 16193 792
rect 16193 758 16201 792
rect 16213 758 16227 792
rect 16227 758 16265 792
rect 16277 758 16299 792
rect 16299 758 16329 792
rect 16341 758 16371 792
rect 16371 758 16393 792
rect 15957 749 16009 758
rect 16021 749 16073 758
rect 16085 749 16137 758
rect 16149 749 16201 758
rect 16213 749 16265 758
rect 16277 749 16329 758
rect 16341 749 16393 758
rect 16405 792 16457 801
rect 16405 758 16409 792
rect 16409 758 16443 792
rect 16443 758 16457 792
rect 16405 749 16457 758
rect 16469 792 16521 801
rect 16469 758 16481 792
rect 16481 758 16515 792
rect 16515 758 16521 792
rect 16469 749 16521 758
rect 16533 792 16585 801
rect 16597 792 16649 801
rect 16661 792 16713 801
rect 16725 792 16777 801
rect 16789 792 16841 801
rect 16853 792 16905 801
rect 16917 792 16969 801
rect 16533 758 16553 792
rect 16553 758 16585 792
rect 16597 758 16625 792
rect 16625 758 16649 792
rect 16661 758 16697 792
rect 16697 758 16713 792
rect 16725 758 16731 792
rect 16731 758 16769 792
rect 16769 758 16777 792
rect 16789 758 16803 792
rect 16803 758 16841 792
rect 16853 758 16875 792
rect 16875 758 16905 792
rect 16917 758 16947 792
rect 16947 758 16969 792
rect 16533 749 16585 758
rect 16597 749 16649 758
rect 16661 749 16713 758
rect 16725 749 16777 758
rect 16789 749 16841 758
rect 16853 749 16905 758
rect 16917 749 16969 758
rect 16981 792 17033 801
rect 16981 758 16985 792
rect 16985 758 17019 792
rect 17019 758 17033 792
rect 16981 749 17033 758
rect 17045 792 17097 801
rect 17045 758 17057 792
rect 17057 758 17091 792
rect 17091 758 17097 792
rect 17045 749 17097 758
rect 17109 792 17161 801
rect 17173 792 17225 801
rect 17237 792 17289 801
rect 17301 792 17353 801
rect 17365 792 17417 801
rect 17429 792 17481 801
rect 17493 792 17545 801
rect 17109 758 17129 792
rect 17129 758 17161 792
rect 17173 758 17201 792
rect 17201 758 17225 792
rect 17237 758 17273 792
rect 17273 758 17289 792
rect 17301 758 17307 792
rect 17307 758 17345 792
rect 17345 758 17353 792
rect 17365 758 17379 792
rect 17379 758 17417 792
rect 17429 758 17451 792
rect 17451 758 17481 792
rect 17493 758 17523 792
rect 17523 758 17545 792
rect 17109 749 17161 758
rect 17173 749 17225 758
rect 17237 749 17289 758
rect 17301 749 17353 758
rect 17365 749 17417 758
rect 17429 749 17481 758
rect 17493 749 17545 758
rect 17557 792 17609 801
rect 17557 758 17561 792
rect 17561 758 17595 792
rect 17595 758 17609 792
rect 17557 749 17609 758
rect 17621 792 17673 801
rect 17621 758 17633 792
rect 17633 758 17667 792
rect 17667 758 17673 792
rect 17621 749 17673 758
rect 17685 792 17737 801
rect 17749 792 17801 801
rect 17813 792 17865 801
rect 17877 792 17929 801
rect 17941 792 17993 801
rect 18005 792 18057 801
rect 18069 792 18121 801
rect 17685 758 17705 792
rect 17705 758 17737 792
rect 17749 758 17777 792
rect 17777 758 17801 792
rect 17813 758 17849 792
rect 17849 758 17865 792
rect 17877 758 17883 792
rect 17883 758 17921 792
rect 17921 758 17929 792
rect 17941 758 17955 792
rect 17955 758 17993 792
rect 18005 758 18027 792
rect 18027 758 18057 792
rect 18069 758 18099 792
rect 18099 758 18121 792
rect 17685 749 17737 758
rect 17749 749 17801 758
rect 17813 749 17865 758
rect 17877 749 17929 758
rect 17941 749 17993 758
rect 18005 749 18057 758
rect 18069 749 18121 758
rect 18133 792 18185 801
rect 18133 758 18137 792
rect 18137 758 18171 792
rect 18171 758 18185 792
rect 18133 749 18185 758
rect 18197 792 18249 801
rect 18197 758 18209 792
rect 18209 758 18243 792
rect 18243 758 18249 792
rect 18197 749 18249 758
rect 18261 792 18313 801
rect 18325 792 18377 801
rect 18389 792 18441 801
rect 18453 792 18505 801
rect 18517 792 18569 801
rect 18581 792 18633 801
rect 18645 792 18697 801
rect 18261 758 18281 792
rect 18281 758 18313 792
rect 18325 758 18353 792
rect 18353 758 18377 792
rect 18389 758 18425 792
rect 18425 758 18441 792
rect 18453 758 18459 792
rect 18459 758 18497 792
rect 18497 758 18505 792
rect 18517 758 18531 792
rect 18531 758 18569 792
rect 18581 758 18603 792
rect 18603 758 18633 792
rect 18645 758 18675 792
rect 18675 758 18697 792
rect 18261 749 18313 758
rect 18325 749 18377 758
rect 18389 749 18441 758
rect 18453 749 18505 758
rect 18517 749 18569 758
rect 18581 749 18633 758
rect 18645 749 18697 758
rect 18709 792 18761 801
rect 18709 758 18713 792
rect 18713 758 18747 792
rect 18747 758 18761 792
rect 18709 749 18761 758
rect 18773 792 18825 801
rect 18773 758 18785 792
rect 18785 758 18819 792
rect 18819 758 18825 792
rect 18773 749 18825 758
rect 18837 749 18889 801
rect 18901 749 18953 801
rect 18965 792 19017 801
rect 18965 758 18983 792
rect 18983 758 19017 792
rect 18965 749 19017 758
rect 19029 792 19081 801
rect 19093 792 19145 801
rect 19157 792 19209 801
rect 19221 792 19273 801
rect 19285 792 19337 801
rect 19349 792 19401 801
rect 19029 758 19055 792
rect 19055 758 19081 792
rect 19093 758 19127 792
rect 19127 758 19145 792
rect 19157 758 19161 792
rect 19161 758 19199 792
rect 19199 758 19209 792
rect 19221 758 19233 792
rect 19233 758 19271 792
rect 19271 758 19273 792
rect 19285 758 19305 792
rect 19305 758 19337 792
rect 19349 758 19377 792
rect 19377 758 19401 792
rect 19029 749 19081 758
rect 19093 749 19145 758
rect 19157 749 19209 758
rect 19221 749 19273 758
rect 19285 749 19337 758
rect 19349 749 19401 758
rect 19413 792 19465 801
rect 19413 758 19415 792
rect 19415 758 19449 792
rect 19449 758 19465 792
rect 19413 749 19465 758
rect 19477 792 19529 801
rect 19477 758 19487 792
rect 19487 758 19521 792
rect 19521 758 19529 792
rect 19477 749 19529 758
rect 19541 792 19593 801
rect 19541 758 19559 792
rect 19559 758 19593 792
rect 19541 749 19593 758
rect 19605 792 19657 801
rect 19669 792 19721 801
rect 19733 792 19785 801
rect 19797 792 19849 801
rect 19861 792 19913 801
rect 19925 792 19977 801
rect 19605 758 19631 792
rect 19631 758 19657 792
rect 19669 758 19703 792
rect 19703 758 19721 792
rect 19733 758 19737 792
rect 19737 758 19775 792
rect 19775 758 19785 792
rect 19797 758 19809 792
rect 19809 758 19847 792
rect 19847 758 19849 792
rect 19861 758 19881 792
rect 19881 758 19913 792
rect 19925 758 19953 792
rect 19953 758 19977 792
rect 19605 749 19657 758
rect 19669 749 19721 758
rect 19733 749 19785 758
rect 19797 749 19849 758
rect 19861 749 19913 758
rect 19925 749 19977 758
rect 19989 792 20041 801
rect 19989 758 19991 792
rect 19991 758 20025 792
rect 20025 758 20041 792
rect 19989 749 20041 758
rect 20053 792 20105 801
rect 20053 758 20063 792
rect 20063 758 20097 792
rect 20097 758 20105 792
rect 20053 749 20105 758
rect 20117 792 20169 801
rect 20117 758 20135 792
rect 20135 758 20169 792
rect 20117 749 20169 758
rect 20181 792 20233 801
rect 20245 792 20297 801
rect 20309 792 20361 801
rect 20373 792 20425 801
rect 20437 792 20489 801
rect 20501 792 20553 801
rect 20181 758 20207 792
rect 20207 758 20233 792
rect 20245 758 20279 792
rect 20279 758 20297 792
rect 20309 758 20313 792
rect 20313 758 20351 792
rect 20351 758 20361 792
rect 20373 758 20385 792
rect 20385 758 20423 792
rect 20423 758 20425 792
rect 20437 758 20457 792
rect 20457 758 20489 792
rect 20501 758 20529 792
rect 20529 758 20553 792
rect 20181 749 20233 758
rect 20245 749 20297 758
rect 20309 749 20361 758
rect 20373 749 20425 758
rect 20437 749 20489 758
rect 20501 749 20553 758
rect 20565 792 20617 801
rect 20565 758 20567 792
rect 20567 758 20601 792
rect 20601 758 20617 792
rect 20565 749 20617 758
rect 20629 792 20681 801
rect 20629 758 20639 792
rect 20639 758 20673 792
rect 20673 758 20681 792
rect 20629 749 20681 758
rect 20693 792 20745 801
rect 20693 758 20711 792
rect 20711 758 20745 792
rect 20693 749 20745 758
rect 20757 792 20809 801
rect 20821 792 20873 801
rect 20885 792 20937 801
rect 20949 792 21001 801
rect 21013 792 21065 801
rect 21077 792 21129 801
rect 20757 758 20783 792
rect 20783 758 20809 792
rect 20821 758 20855 792
rect 20855 758 20873 792
rect 20885 758 20889 792
rect 20889 758 20927 792
rect 20927 758 20937 792
rect 20949 758 20961 792
rect 20961 758 20999 792
rect 20999 758 21001 792
rect 21013 758 21033 792
rect 21033 758 21065 792
rect 21077 758 21105 792
rect 21105 758 21129 792
rect 20757 749 20809 758
rect 20821 749 20873 758
rect 20885 749 20937 758
rect 20949 749 21001 758
rect 21013 749 21065 758
rect 21077 749 21129 758
rect 21141 792 21193 801
rect 21141 758 21143 792
rect 21143 758 21177 792
rect 21177 758 21193 792
rect 21141 749 21193 758
rect 21205 792 21257 801
rect 21205 758 21215 792
rect 21215 758 21249 792
rect 21249 758 21257 792
rect 21205 749 21257 758
rect 21269 792 21321 801
rect 21269 758 21287 792
rect 21287 758 21321 792
rect 21269 749 21321 758
rect 21333 792 21385 801
rect 21397 792 21449 801
rect 21461 792 21513 801
rect 21525 792 21577 801
rect 21589 792 21641 801
rect 21653 792 21705 801
rect 21333 758 21359 792
rect 21359 758 21385 792
rect 21397 758 21431 792
rect 21431 758 21449 792
rect 21461 758 21465 792
rect 21465 758 21503 792
rect 21503 758 21513 792
rect 21525 758 21537 792
rect 21537 758 21575 792
rect 21575 758 21577 792
rect 21589 758 21609 792
rect 21609 758 21641 792
rect 21653 758 21681 792
rect 21681 758 21705 792
rect 21333 749 21385 758
rect 21397 749 21449 758
rect 21461 749 21513 758
rect 21525 749 21577 758
rect 21589 749 21641 758
rect 21653 749 21705 758
rect 21717 792 21769 801
rect 21717 758 21719 792
rect 21719 758 21753 792
rect 21753 758 21769 792
rect 21717 749 21769 758
rect 21781 792 21833 801
rect 21781 758 21791 792
rect 21791 758 21825 792
rect 21825 758 21833 792
rect 21781 749 21833 758
rect 21845 792 21897 801
rect 21845 758 21863 792
rect 21863 758 21897 792
rect 21845 749 21897 758
rect 21909 792 21961 801
rect 21909 758 21935 792
rect 21935 758 21961 792
rect 21909 749 21961 758
rect 22236 785 22288 802
rect 22236 760 22288 772
rect 22236 726 22248 760
rect 22248 726 22282 760
rect 22282 726 22288 760
rect 22236 720 22288 726
rect 23407 702 23459 711
rect 23478 702 23530 711
rect 23549 702 23601 711
rect 23620 702 23672 711
rect 23691 702 23743 711
rect 23762 702 23814 711
rect 23833 702 23885 711
rect 23904 702 23956 711
rect 23975 702 24027 711
rect 24046 702 24098 711
rect 1545 662 1597 671
rect 1610 662 1662 671
rect 1675 662 1727 671
rect 1740 662 1792 671
rect 1545 628 1557 662
rect 1557 628 1595 662
rect 1595 628 1597 662
rect 1610 628 1629 662
rect 1629 628 1662 662
rect 1675 628 1701 662
rect 1701 628 1727 662
rect 1740 628 1773 662
rect 1773 628 1792 662
rect 1545 619 1597 628
rect 1610 619 1662 628
rect 1675 619 1727 628
rect 1740 619 1792 628
rect 1805 662 1857 671
rect 1805 628 1811 662
rect 1811 628 1845 662
rect 1845 628 1857 662
rect 1805 619 1857 628
rect 1870 662 1922 671
rect 1870 628 1883 662
rect 1883 628 1917 662
rect 1917 628 1922 662
rect 1870 619 1922 628
rect 1935 662 1987 671
rect 2000 662 2052 671
rect 2065 662 2117 671
rect 2130 662 2182 671
rect 2195 662 2247 671
rect 2260 662 2312 671
rect 2325 662 2377 671
rect 2390 662 2442 671
rect 1935 628 1955 662
rect 1955 628 1987 662
rect 2000 628 2027 662
rect 2027 628 2052 662
rect 2065 628 2099 662
rect 2099 628 2117 662
rect 2130 628 2133 662
rect 2133 628 2171 662
rect 2171 628 2182 662
rect 2195 628 2205 662
rect 2205 628 2243 662
rect 2243 628 2247 662
rect 2260 628 2277 662
rect 2277 628 2312 662
rect 2325 628 2349 662
rect 2349 628 2377 662
rect 2390 628 2421 662
rect 2421 628 2442 662
rect 1935 619 1987 628
rect 2000 619 2052 628
rect 2065 619 2117 628
rect 2130 619 2182 628
rect 2195 619 2247 628
rect 2260 619 2312 628
rect 2325 619 2377 628
rect 2390 619 2442 628
rect 2455 662 2507 671
rect 2455 628 2459 662
rect 2459 628 2493 662
rect 2493 628 2507 662
rect 2455 619 2507 628
rect 2520 662 2572 671
rect 2520 628 2531 662
rect 2531 628 2565 662
rect 2565 628 2572 662
rect 2520 619 2572 628
rect 2585 662 2637 671
rect 2585 628 2603 662
rect 2603 628 2637 662
rect 2585 619 2637 628
rect 2650 662 2702 671
rect 2715 662 2767 671
rect 2780 662 2832 671
rect 2845 662 2897 671
rect 2910 662 2962 671
rect 2975 662 3027 671
rect 3040 662 3092 671
rect 2650 628 2675 662
rect 2675 628 2702 662
rect 2715 628 2747 662
rect 2747 628 2767 662
rect 2780 628 2781 662
rect 2781 628 2819 662
rect 2819 628 2832 662
rect 2845 628 2853 662
rect 2853 628 2891 662
rect 2891 628 2897 662
rect 2910 628 2925 662
rect 2925 628 2962 662
rect 2975 628 2997 662
rect 2997 628 3027 662
rect 3040 628 3069 662
rect 3069 628 3092 662
rect 2650 619 2702 628
rect 2715 619 2767 628
rect 2780 619 2832 628
rect 2845 619 2897 628
rect 2910 619 2962 628
rect 2975 619 3027 628
rect 3040 619 3092 628
rect 3105 619 3157 671
rect 3170 619 3222 671
rect 3235 662 3287 671
rect 3235 628 3267 662
rect 3267 628 3287 662
rect 3235 619 3287 628
rect 3300 662 3352 671
rect 3300 628 3305 662
rect 3305 628 3339 662
rect 3339 628 3352 662
rect 3300 619 3352 628
rect 3365 662 3417 671
rect 3365 628 3377 662
rect 3377 628 3411 662
rect 3411 628 3417 662
rect 3365 619 3417 628
rect 3430 662 3482 671
rect 3495 662 3547 671
rect 3560 662 3612 671
rect 3625 662 3677 671
rect 3690 662 3742 671
rect 3755 662 3807 671
rect 3820 662 3872 671
rect 3885 662 3937 671
rect 3430 628 3449 662
rect 3449 628 3482 662
rect 3495 628 3521 662
rect 3521 628 3547 662
rect 3560 628 3593 662
rect 3593 628 3612 662
rect 3625 628 3627 662
rect 3627 628 3665 662
rect 3665 628 3677 662
rect 3690 628 3699 662
rect 3699 628 3737 662
rect 3737 628 3742 662
rect 3755 628 3771 662
rect 3771 628 3807 662
rect 3820 628 3843 662
rect 3843 628 3872 662
rect 3885 628 3915 662
rect 3915 628 3937 662
rect 3430 619 3482 628
rect 3495 619 3547 628
rect 3560 619 3612 628
rect 3625 619 3677 628
rect 3690 619 3742 628
rect 3755 619 3807 628
rect 3820 619 3872 628
rect 3885 619 3937 628
rect 3950 662 4002 671
rect 3950 628 3953 662
rect 3953 628 3987 662
rect 3987 628 4002 662
rect 3950 619 4002 628
rect 4015 662 4067 671
rect 4015 628 4025 662
rect 4025 628 4059 662
rect 4059 628 4067 662
rect 4015 619 4067 628
rect 4080 662 4132 671
rect 4080 628 4097 662
rect 4097 628 4131 662
rect 4131 628 4132 662
rect 4080 619 4132 628
rect 4144 662 4196 671
rect 4208 662 4260 671
rect 4272 662 4324 671
rect 4336 662 4388 671
rect 4400 662 4452 671
rect 4464 662 4516 671
rect 4144 628 4169 662
rect 4169 628 4196 662
rect 4208 628 4241 662
rect 4241 628 4260 662
rect 4272 628 4275 662
rect 4275 628 4313 662
rect 4313 628 4324 662
rect 4336 628 4347 662
rect 4347 628 4385 662
rect 4385 628 4388 662
rect 4400 628 4419 662
rect 4419 628 4452 662
rect 4464 628 4491 662
rect 4491 628 4516 662
rect 4144 619 4196 628
rect 4208 619 4260 628
rect 4272 619 4324 628
rect 4336 619 4388 628
rect 4400 619 4452 628
rect 4464 619 4516 628
rect 4528 662 4580 671
rect 4528 628 4529 662
rect 4529 628 4563 662
rect 4563 628 4580 662
rect 4528 619 4580 628
rect 4592 662 4644 671
rect 4592 628 4601 662
rect 4601 628 4635 662
rect 4635 628 4644 662
rect 4592 619 4644 628
rect 4656 662 4708 671
rect 4656 628 4673 662
rect 4673 628 4707 662
rect 4707 628 4708 662
rect 4656 619 4708 628
rect 4720 662 4772 671
rect 4784 662 4836 671
rect 4848 662 4900 671
rect 4912 662 4964 671
rect 4976 662 5028 671
rect 5040 662 5092 671
rect 4720 628 4745 662
rect 4745 628 4772 662
rect 4784 628 4817 662
rect 4817 628 4836 662
rect 4848 628 4851 662
rect 4851 628 4889 662
rect 4889 628 4900 662
rect 4912 628 4923 662
rect 4923 628 4961 662
rect 4961 628 4964 662
rect 4976 628 4995 662
rect 4995 628 5028 662
rect 5040 628 5067 662
rect 5067 628 5092 662
rect 4720 619 4772 628
rect 4784 619 4836 628
rect 4848 619 4900 628
rect 4912 619 4964 628
rect 4976 619 5028 628
rect 5040 619 5092 628
rect 5104 662 5156 671
rect 5104 628 5105 662
rect 5105 628 5139 662
rect 5139 628 5156 662
rect 5104 619 5156 628
rect 5168 662 5220 671
rect 5168 628 5177 662
rect 5177 628 5211 662
rect 5211 628 5220 662
rect 5168 619 5220 628
rect 5232 662 5284 671
rect 5232 628 5249 662
rect 5249 628 5283 662
rect 5283 628 5284 662
rect 5232 619 5284 628
rect 5296 662 5348 671
rect 5360 662 5412 671
rect 5424 662 5476 671
rect 5488 662 5540 671
rect 5552 662 5604 671
rect 5616 662 5668 671
rect 5296 628 5321 662
rect 5321 628 5348 662
rect 5360 628 5393 662
rect 5393 628 5412 662
rect 5424 628 5427 662
rect 5427 628 5465 662
rect 5465 628 5476 662
rect 5488 628 5499 662
rect 5499 628 5537 662
rect 5537 628 5540 662
rect 5552 628 5571 662
rect 5571 628 5604 662
rect 5616 628 5643 662
rect 5643 628 5668 662
rect 5296 619 5348 628
rect 5360 619 5412 628
rect 5424 619 5476 628
rect 5488 619 5540 628
rect 5552 619 5604 628
rect 5616 619 5668 628
rect 5680 662 5732 671
rect 5680 628 5681 662
rect 5681 628 5715 662
rect 5715 628 5732 662
rect 5680 619 5732 628
rect 5744 662 5796 671
rect 5744 628 5753 662
rect 5753 628 5787 662
rect 5787 628 5796 662
rect 5744 619 5796 628
rect 5808 662 5860 671
rect 5808 628 5825 662
rect 5825 628 5859 662
rect 5859 628 5860 662
rect 5808 619 5860 628
rect 5872 662 5924 671
rect 5936 662 5988 671
rect 6000 662 6052 671
rect 6064 662 6116 671
rect 23407 668 23408 702
rect 23408 668 23446 702
rect 23446 668 23459 702
rect 23478 668 23480 702
rect 23480 668 23518 702
rect 23518 668 23530 702
rect 23549 668 23552 702
rect 23552 668 23590 702
rect 23590 668 23601 702
rect 23620 668 23624 702
rect 23624 668 23662 702
rect 23662 668 23672 702
rect 23691 668 23696 702
rect 23696 668 23734 702
rect 23734 668 23743 702
rect 23762 668 23768 702
rect 23768 668 23806 702
rect 23806 668 23814 702
rect 23833 668 23840 702
rect 23840 668 23878 702
rect 23878 668 23885 702
rect 23904 668 23912 702
rect 23912 668 23950 702
rect 23950 668 23956 702
rect 23975 668 23984 702
rect 23984 668 24022 702
rect 24022 668 24027 702
rect 24046 668 24056 702
rect 24056 668 24094 702
rect 24094 668 24098 702
rect 5872 628 5897 662
rect 5897 628 5924 662
rect 5936 628 5969 662
rect 5969 628 5988 662
rect 6000 628 6003 662
rect 6003 628 6041 662
rect 6041 628 6052 662
rect 6064 628 6075 662
rect 6075 628 6113 662
rect 6113 628 6116 662
rect 23407 659 23459 668
rect 23478 659 23530 668
rect 23549 659 23601 668
rect 23620 659 23672 668
rect 23691 659 23743 668
rect 23762 659 23814 668
rect 23833 659 23885 668
rect 23904 659 23956 668
rect 23975 659 24027 668
rect 24046 659 24098 668
rect 5872 619 5924 628
rect 5936 619 5988 628
rect 6000 619 6052 628
rect 6064 619 6116 628
rect 7616 636 7668 645
rect 7681 636 7733 645
rect 7616 602 7641 636
rect 7641 602 7668 636
rect 7681 602 7713 636
rect 7713 602 7733 636
rect 7616 593 7668 602
rect 7681 593 7733 602
rect 7746 636 7798 645
rect 7746 602 7751 636
rect 7751 602 7785 636
rect 7785 602 7798 636
rect 7746 593 7798 602
rect 7811 636 7863 645
rect 7811 602 7823 636
rect 7823 602 7857 636
rect 7857 602 7863 636
rect 7811 593 7863 602
rect 7876 636 7928 645
rect 7941 636 7993 645
rect 8006 636 8058 645
rect 8071 636 8123 645
rect 8136 636 8188 645
rect 8201 636 8253 645
rect 8266 636 8318 645
rect 8331 636 8383 645
rect 7876 602 7895 636
rect 7895 602 7928 636
rect 7941 602 7967 636
rect 7967 602 7993 636
rect 8006 602 8039 636
rect 8039 602 8058 636
rect 8071 602 8073 636
rect 8073 602 8111 636
rect 8111 602 8123 636
rect 8136 602 8145 636
rect 8145 602 8183 636
rect 8183 602 8188 636
rect 8201 602 8217 636
rect 8217 602 8253 636
rect 8266 602 8289 636
rect 8289 602 8318 636
rect 8331 602 8361 636
rect 8361 602 8383 636
rect 7876 593 7928 602
rect 7941 593 7993 602
rect 8006 593 8058 602
rect 8071 593 8123 602
rect 8136 593 8188 602
rect 8201 593 8253 602
rect 8266 593 8318 602
rect 8331 593 8383 602
rect 8396 636 8448 645
rect 8396 602 8399 636
rect 8399 602 8433 636
rect 8433 602 8448 636
rect 8396 593 8448 602
rect 8461 636 8513 645
rect 8461 602 8471 636
rect 8471 602 8505 636
rect 8505 602 8513 636
rect 8461 593 8513 602
rect 8526 636 8578 645
rect 8526 602 8543 636
rect 8543 602 8577 636
rect 8577 602 8578 636
rect 8526 593 8578 602
rect 8591 636 8643 645
rect 8656 636 8708 645
rect 8721 636 8773 645
rect 8786 636 8838 645
rect 8851 636 8903 645
rect 8916 636 8968 645
rect 8981 636 9033 645
rect 8591 602 8615 636
rect 8615 602 8643 636
rect 8656 602 8687 636
rect 8687 602 8708 636
rect 8721 602 8759 636
rect 8759 602 8773 636
rect 8786 602 8793 636
rect 8793 602 8831 636
rect 8831 602 8838 636
rect 8851 602 8865 636
rect 8865 602 8903 636
rect 8916 602 8937 636
rect 8937 602 8968 636
rect 8981 602 9009 636
rect 9009 602 9033 636
rect 8591 593 8643 602
rect 8656 593 8708 602
rect 8721 593 8773 602
rect 8786 593 8838 602
rect 8851 593 8903 602
rect 8916 593 8968 602
rect 8981 593 9033 602
rect 9046 636 9098 645
rect 9046 602 9047 636
rect 9047 602 9081 636
rect 9081 602 9098 636
rect 9046 593 9098 602
rect 9111 636 9163 645
rect 9111 602 9119 636
rect 9119 602 9153 636
rect 9153 602 9163 636
rect 9111 593 9163 602
rect 9176 636 9228 645
rect 9176 602 9191 636
rect 9191 602 9225 636
rect 9225 602 9228 636
rect 9176 593 9228 602
rect 9241 636 9293 645
rect 9306 636 9358 645
rect 9241 602 9263 636
rect 9263 602 9293 636
rect 9306 602 9335 636
rect 9335 602 9358 636
rect 9241 593 9293 602
rect 9306 593 9358 602
rect 9371 593 9423 645
rect 9436 593 9488 645
rect 9501 636 9553 645
rect 9566 636 9618 645
rect 9631 636 9683 645
rect 9696 636 9748 645
rect 9761 636 9813 645
rect 9826 636 9878 645
rect 9501 602 9533 636
rect 9533 602 9553 636
rect 9566 602 9567 636
rect 9567 602 9605 636
rect 9605 602 9618 636
rect 9631 602 9639 636
rect 9639 602 9677 636
rect 9677 602 9683 636
rect 9696 602 9711 636
rect 9711 602 9748 636
rect 9761 602 9783 636
rect 9783 602 9813 636
rect 9826 602 9855 636
rect 9855 602 9878 636
rect 9501 593 9553 602
rect 9566 593 9618 602
rect 9631 593 9683 602
rect 9696 593 9748 602
rect 9761 593 9813 602
rect 9826 593 9878 602
rect 9891 636 9943 645
rect 9891 602 9893 636
rect 9893 602 9927 636
rect 9927 602 9943 636
rect 9891 593 9943 602
rect 9956 636 10008 645
rect 9956 602 9965 636
rect 9965 602 9999 636
rect 9999 602 10008 636
rect 9956 593 10008 602
rect 10021 636 10073 645
rect 10021 602 10037 636
rect 10037 602 10071 636
rect 10071 602 10073 636
rect 10021 593 10073 602
rect 10086 636 10138 645
rect 10151 636 10203 645
rect 10216 636 10268 645
rect 10281 636 10333 645
rect 10346 636 10398 645
rect 10411 636 10463 645
rect 10476 636 10528 645
rect 10086 602 10109 636
rect 10109 602 10138 636
rect 10151 602 10181 636
rect 10181 602 10203 636
rect 10216 602 10253 636
rect 10253 602 10268 636
rect 10281 602 10287 636
rect 10287 602 10325 636
rect 10325 602 10333 636
rect 10346 602 10359 636
rect 10359 602 10397 636
rect 10397 602 10398 636
rect 10411 602 10431 636
rect 10431 602 10463 636
rect 10476 602 10503 636
rect 10503 602 10528 636
rect 10086 593 10138 602
rect 10151 593 10203 602
rect 10216 593 10268 602
rect 10281 593 10333 602
rect 10346 593 10398 602
rect 10411 593 10463 602
rect 10476 593 10528 602
rect 10541 636 10593 645
rect 10541 602 10575 636
rect 10575 602 10593 636
rect 10541 593 10593 602
rect 10606 636 10658 645
rect 10606 602 10613 636
rect 10613 602 10647 636
rect 10647 602 10658 636
rect 10606 593 10658 602
rect 10671 636 10723 645
rect 10671 602 10685 636
rect 10685 602 10719 636
rect 10719 602 10723 636
rect 10671 593 10723 602
rect 10736 636 10788 645
rect 10800 636 10852 645
rect 10864 636 10916 645
rect 10928 636 10980 645
rect 10992 636 11044 645
rect 11056 636 11108 645
rect 11120 636 11172 645
rect 10736 602 10757 636
rect 10757 602 10788 636
rect 10800 602 10829 636
rect 10829 602 10852 636
rect 10864 602 10901 636
rect 10901 602 10916 636
rect 10928 602 10935 636
rect 10935 602 10973 636
rect 10973 602 10980 636
rect 10992 602 11007 636
rect 11007 602 11044 636
rect 11056 602 11079 636
rect 11079 602 11108 636
rect 11120 602 11151 636
rect 11151 602 11172 636
rect 10736 593 10788 602
rect 10800 593 10852 602
rect 10864 593 10916 602
rect 10928 593 10980 602
rect 10992 593 11044 602
rect 11056 593 11108 602
rect 11120 593 11172 602
rect 11184 636 11236 645
rect 11184 602 11189 636
rect 11189 602 11223 636
rect 11223 602 11236 636
rect 11184 593 11236 602
rect 11248 636 11300 645
rect 11248 602 11261 636
rect 11261 602 11295 636
rect 11295 602 11300 636
rect 11248 593 11300 602
rect 11312 636 11364 645
rect 11376 636 11428 645
rect 11440 636 11492 645
rect 11504 636 11556 645
rect 11568 636 11620 645
rect 11632 636 11684 645
rect 11696 636 11748 645
rect 11312 602 11333 636
rect 11333 602 11364 636
rect 11376 602 11405 636
rect 11405 602 11428 636
rect 11440 602 11477 636
rect 11477 602 11492 636
rect 11504 602 11511 636
rect 11511 602 11549 636
rect 11549 602 11556 636
rect 11568 602 11583 636
rect 11583 602 11620 636
rect 11632 602 11655 636
rect 11655 602 11684 636
rect 11696 602 11727 636
rect 11727 602 11748 636
rect 11312 593 11364 602
rect 11376 593 11428 602
rect 11440 593 11492 602
rect 11504 593 11556 602
rect 11568 593 11620 602
rect 11632 593 11684 602
rect 11696 593 11748 602
rect 11760 636 11812 645
rect 11760 602 11765 636
rect 11765 602 11799 636
rect 11799 602 11812 636
rect 11760 593 11812 602
rect 11824 636 11876 645
rect 12022 636 12074 645
rect 12087 636 12139 645
rect 12152 636 12204 645
rect 12217 636 12269 645
rect 12282 636 12334 645
rect 12347 636 12399 645
rect 11824 602 11837 636
rect 11837 602 11871 636
rect 11871 602 11876 636
rect 12022 602 12053 636
rect 12053 602 12074 636
rect 12087 602 12125 636
rect 12125 602 12139 636
rect 12152 602 12159 636
rect 12159 602 12197 636
rect 12197 602 12204 636
rect 12217 602 12231 636
rect 12231 602 12269 636
rect 12282 602 12303 636
rect 12303 602 12334 636
rect 12347 602 12375 636
rect 12375 602 12399 636
rect 11824 593 11876 602
rect 12022 593 12074 602
rect 12087 593 12139 602
rect 12152 593 12204 602
rect 12217 593 12269 602
rect 12282 593 12334 602
rect 12347 593 12399 602
rect 12412 636 12464 645
rect 12412 602 12413 636
rect 12413 602 12447 636
rect 12447 602 12464 636
rect 12412 593 12464 602
rect 12477 636 12529 645
rect 12477 602 12485 636
rect 12485 602 12519 636
rect 12519 602 12529 636
rect 12477 593 12529 602
rect 12542 593 12594 645
rect 12607 593 12659 645
rect 12672 636 12724 645
rect 12672 602 12683 636
rect 12683 602 12717 636
rect 12717 602 12724 636
rect 12672 593 12724 602
rect 12737 636 12789 645
rect 12737 602 12755 636
rect 12755 602 12789 636
rect 12737 593 12789 602
rect 12802 636 12854 645
rect 12867 636 12919 645
rect 12932 636 12984 645
rect 12997 636 13049 645
rect 13062 636 13114 645
rect 13127 636 13179 645
rect 13192 636 13244 645
rect 12802 602 12827 636
rect 12827 602 12854 636
rect 12867 602 12899 636
rect 12899 602 12919 636
rect 12932 602 12933 636
rect 12933 602 12971 636
rect 12971 602 12984 636
rect 12997 602 13005 636
rect 13005 602 13043 636
rect 13043 602 13049 636
rect 13062 602 13077 636
rect 13077 602 13114 636
rect 13127 602 13149 636
rect 13149 602 13179 636
rect 13192 602 13221 636
rect 13221 602 13244 636
rect 12802 593 12854 602
rect 12867 593 12919 602
rect 12932 593 12984 602
rect 12997 593 13049 602
rect 13062 593 13114 602
rect 13127 593 13179 602
rect 13192 593 13244 602
rect 13257 636 13309 645
rect 13257 602 13259 636
rect 13259 602 13293 636
rect 13293 602 13309 636
rect 13257 593 13309 602
rect 13322 636 13374 645
rect 13322 602 13331 636
rect 13331 602 13365 636
rect 13365 602 13374 636
rect 13322 593 13374 602
rect 13387 636 13439 645
rect 13387 602 13403 636
rect 13403 602 13437 636
rect 13437 602 13439 636
rect 13387 593 13439 602
rect 13452 636 13504 645
rect 13517 636 13569 645
rect 13582 636 13634 645
rect 13647 636 13699 645
rect 13712 636 13764 645
rect 13777 636 13829 645
rect 13842 636 13894 645
rect 13452 602 13475 636
rect 13475 602 13504 636
rect 13517 602 13547 636
rect 13547 602 13569 636
rect 13582 602 13619 636
rect 13619 602 13634 636
rect 13647 602 13653 636
rect 13653 602 13691 636
rect 13691 602 13699 636
rect 13712 602 13725 636
rect 13725 602 13763 636
rect 13763 602 13764 636
rect 13777 602 13797 636
rect 13797 602 13829 636
rect 13842 602 13869 636
rect 13869 602 13894 636
rect 13452 593 13504 602
rect 13517 593 13569 602
rect 13582 593 13634 602
rect 13647 593 13699 602
rect 13712 593 13764 602
rect 13777 593 13829 602
rect 13842 593 13894 602
rect 13907 636 13959 645
rect 13907 602 13941 636
rect 13941 602 13959 636
rect 13907 593 13959 602
rect 13972 636 14024 645
rect 13972 602 13979 636
rect 13979 602 14013 636
rect 14013 602 14024 636
rect 13972 593 14024 602
rect 14037 636 14089 645
rect 14037 602 14051 636
rect 14051 602 14085 636
rect 14085 602 14089 636
rect 14037 593 14089 602
rect 14102 636 14154 645
rect 14167 636 14219 645
rect 14232 636 14284 645
rect 14297 636 14349 645
rect 14362 636 14414 645
rect 14427 636 14479 645
rect 14492 636 14544 645
rect 14557 636 14609 645
rect 14102 602 14123 636
rect 14123 602 14154 636
rect 14167 602 14195 636
rect 14195 602 14219 636
rect 14232 602 14267 636
rect 14267 602 14284 636
rect 14297 602 14301 636
rect 14301 602 14339 636
rect 14339 602 14349 636
rect 14362 602 14373 636
rect 14373 602 14411 636
rect 14411 602 14414 636
rect 14427 602 14445 636
rect 14445 602 14479 636
rect 14492 602 14517 636
rect 14517 602 14544 636
rect 14557 602 14589 636
rect 14589 602 14609 636
rect 14102 593 14154 602
rect 14167 593 14219 602
rect 14232 593 14284 602
rect 14297 593 14349 602
rect 14362 593 14414 602
rect 14427 593 14479 602
rect 14492 593 14544 602
rect 14557 593 14609 602
rect 14622 636 14674 645
rect 14622 602 14627 636
rect 14627 602 14661 636
rect 14661 602 14674 636
rect 14622 593 14674 602
rect 14687 636 14739 645
rect 14687 602 14699 636
rect 14699 602 14733 636
rect 14733 602 14739 636
rect 14687 593 14739 602
rect 14752 636 14804 645
rect 14817 636 14869 645
rect 14882 636 14934 645
rect 14947 636 14999 645
rect 15012 636 15064 645
rect 15077 636 15129 645
rect 15142 636 15194 645
rect 15206 636 15258 645
rect 14752 602 14771 636
rect 14771 602 14804 636
rect 14817 602 14843 636
rect 14843 602 14869 636
rect 14882 602 14915 636
rect 14915 602 14934 636
rect 14947 602 14949 636
rect 14949 602 14987 636
rect 14987 602 14999 636
rect 15012 602 15021 636
rect 15021 602 15059 636
rect 15059 602 15064 636
rect 15077 602 15093 636
rect 15093 602 15129 636
rect 15142 602 15165 636
rect 15165 602 15194 636
rect 15206 602 15237 636
rect 15237 602 15258 636
rect 14752 593 14804 602
rect 14817 593 14869 602
rect 14882 593 14934 602
rect 14947 593 14999 602
rect 15012 593 15064 602
rect 15077 593 15129 602
rect 15142 593 15194 602
rect 15206 593 15258 602
rect 15270 636 15322 645
rect 15270 602 15275 636
rect 15275 602 15309 636
rect 15309 602 15322 636
rect 15270 593 15322 602
rect 15334 636 15386 645
rect 15334 602 15347 636
rect 15347 602 15381 636
rect 15381 602 15386 636
rect 15334 593 15386 602
rect 15398 636 15450 645
rect 15462 636 15514 645
rect 15526 636 15578 645
rect 15590 636 15642 645
rect 15654 636 15706 645
rect 15398 602 15419 636
rect 15419 602 15450 636
rect 15462 602 15491 636
rect 15491 602 15514 636
rect 15526 602 15563 636
rect 15563 602 15578 636
rect 15590 602 15597 636
rect 15597 602 15635 636
rect 15635 602 15642 636
rect 15654 602 15669 636
rect 15669 602 15706 636
rect 15398 593 15450 602
rect 15462 593 15514 602
rect 15526 593 15578 602
rect 15590 593 15642 602
rect 15654 593 15706 602
rect 15718 593 15770 645
rect 15782 636 15834 645
rect 15846 636 15898 645
rect 15910 636 15962 645
rect 15782 602 15833 636
rect 15833 602 15834 636
rect 15846 602 15867 636
rect 15867 602 15898 636
rect 15910 602 15939 636
rect 15939 602 15962 636
rect 15782 593 15834 602
rect 15846 593 15898 602
rect 15910 593 15962 602
rect 15974 636 16026 645
rect 15974 602 15977 636
rect 15977 602 16011 636
rect 16011 602 16026 636
rect 15974 593 16026 602
rect 16038 636 16090 645
rect 16038 602 16049 636
rect 16049 602 16083 636
rect 16083 602 16090 636
rect 16038 593 16090 602
rect 16102 636 16154 645
rect 16166 636 16218 645
rect 16230 636 16282 645
rect 16294 636 16346 645
rect 16358 636 16410 645
rect 16422 636 16474 645
rect 16486 636 16538 645
rect 16102 602 16121 636
rect 16121 602 16154 636
rect 16166 602 16193 636
rect 16193 602 16218 636
rect 16230 602 16265 636
rect 16265 602 16282 636
rect 16294 602 16299 636
rect 16299 602 16337 636
rect 16337 602 16346 636
rect 16358 602 16371 636
rect 16371 602 16409 636
rect 16409 602 16410 636
rect 16422 602 16443 636
rect 16443 602 16474 636
rect 16486 602 16515 636
rect 16515 602 16538 636
rect 16102 593 16154 602
rect 16166 593 16218 602
rect 16230 593 16282 602
rect 16294 593 16346 602
rect 16358 593 16410 602
rect 16422 593 16474 602
rect 16486 593 16538 602
rect 16550 636 16602 645
rect 16550 602 16553 636
rect 16553 602 16587 636
rect 16587 602 16602 636
rect 16550 593 16602 602
rect 16614 636 16666 645
rect 16614 602 16625 636
rect 16625 602 16659 636
rect 16659 602 16666 636
rect 16614 593 16666 602
rect 16678 636 16730 645
rect 16742 636 16794 645
rect 16806 636 16858 645
rect 16870 636 16922 645
rect 16934 636 16986 645
rect 16998 636 17050 645
rect 17062 636 17114 645
rect 16678 602 16697 636
rect 16697 602 16730 636
rect 16742 602 16769 636
rect 16769 602 16794 636
rect 16806 602 16841 636
rect 16841 602 16858 636
rect 16870 602 16875 636
rect 16875 602 16913 636
rect 16913 602 16922 636
rect 16934 602 16947 636
rect 16947 602 16985 636
rect 16985 602 16986 636
rect 16998 602 17019 636
rect 17019 602 17050 636
rect 17062 602 17091 636
rect 17091 602 17114 636
rect 16678 593 16730 602
rect 16742 593 16794 602
rect 16806 593 16858 602
rect 16870 593 16922 602
rect 16934 593 16986 602
rect 16998 593 17050 602
rect 17062 593 17114 602
rect 17126 636 17178 645
rect 17126 602 17129 636
rect 17129 602 17163 636
rect 17163 602 17178 636
rect 17126 593 17178 602
rect 17190 636 17242 645
rect 17190 602 17201 636
rect 17201 602 17235 636
rect 17235 602 17242 636
rect 17190 593 17242 602
rect 17254 636 17306 645
rect 17318 636 17370 645
rect 17382 636 17434 645
rect 17446 636 17498 645
rect 17510 636 17562 645
rect 17574 636 17626 645
rect 17638 636 17690 645
rect 17254 602 17273 636
rect 17273 602 17306 636
rect 17318 602 17345 636
rect 17345 602 17370 636
rect 17382 602 17417 636
rect 17417 602 17434 636
rect 17446 602 17451 636
rect 17451 602 17489 636
rect 17489 602 17498 636
rect 17510 602 17523 636
rect 17523 602 17561 636
rect 17561 602 17562 636
rect 17574 602 17595 636
rect 17595 602 17626 636
rect 17638 602 17667 636
rect 17667 602 17690 636
rect 17254 593 17306 602
rect 17318 593 17370 602
rect 17382 593 17434 602
rect 17446 593 17498 602
rect 17510 593 17562 602
rect 17574 593 17626 602
rect 17638 593 17690 602
rect 17702 636 17754 645
rect 17702 602 17705 636
rect 17705 602 17739 636
rect 17739 602 17754 636
rect 17702 593 17754 602
rect 17766 636 17818 645
rect 17766 602 17777 636
rect 17777 602 17811 636
rect 17811 602 17818 636
rect 17766 593 17818 602
rect 17830 636 17882 645
rect 17894 636 17946 645
rect 17958 636 18010 645
rect 18022 636 18074 645
rect 18086 636 18138 645
rect 18150 636 18202 645
rect 18214 636 18266 645
rect 17830 602 17849 636
rect 17849 602 17882 636
rect 17894 602 17921 636
rect 17921 602 17946 636
rect 17958 602 17993 636
rect 17993 602 18010 636
rect 18022 602 18027 636
rect 18027 602 18065 636
rect 18065 602 18074 636
rect 18086 602 18099 636
rect 18099 602 18137 636
rect 18137 602 18138 636
rect 18150 602 18171 636
rect 18171 602 18202 636
rect 18214 602 18243 636
rect 18243 602 18266 636
rect 17830 593 17882 602
rect 17894 593 17946 602
rect 17958 593 18010 602
rect 18022 593 18074 602
rect 18086 593 18138 602
rect 18150 593 18202 602
rect 18214 593 18266 602
rect 18278 636 18330 645
rect 18278 602 18281 636
rect 18281 602 18315 636
rect 18315 602 18330 636
rect 18278 593 18330 602
rect 18342 636 18394 645
rect 18342 602 18353 636
rect 18353 602 18387 636
rect 18387 602 18394 636
rect 18342 593 18394 602
rect 18406 636 18458 645
rect 18470 636 18522 645
rect 18534 636 18586 645
rect 18598 636 18650 645
rect 18662 636 18714 645
rect 18726 636 18778 645
rect 18790 636 18842 645
rect 18406 602 18425 636
rect 18425 602 18458 636
rect 18470 602 18497 636
rect 18497 602 18522 636
rect 18534 602 18569 636
rect 18569 602 18586 636
rect 18598 602 18603 636
rect 18603 602 18641 636
rect 18641 602 18650 636
rect 18662 602 18675 636
rect 18675 602 18713 636
rect 18713 602 18714 636
rect 18726 602 18747 636
rect 18747 602 18778 636
rect 18790 602 18819 636
rect 18819 602 18842 636
rect 18406 593 18458 602
rect 18470 593 18522 602
rect 18534 593 18586 602
rect 18598 593 18650 602
rect 18662 593 18714 602
rect 18726 593 18778 602
rect 18790 593 18842 602
rect 18854 593 18906 645
rect 18918 593 18970 645
rect 18982 636 19034 645
rect 18982 602 18983 636
rect 18983 602 19017 636
rect 19017 602 19034 636
rect 18982 593 19034 602
rect 19046 636 19098 645
rect 19046 602 19055 636
rect 19055 602 19089 636
rect 19089 602 19098 636
rect 19046 593 19098 602
rect 19110 636 19162 645
rect 19110 602 19127 636
rect 19127 602 19161 636
rect 19161 602 19162 636
rect 19110 593 19162 602
rect 19174 636 19226 645
rect 19238 636 19290 645
rect 19302 636 19354 645
rect 19366 636 19418 645
rect 19430 636 19482 645
rect 19494 636 19546 645
rect 19174 602 19199 636
rect 19199 602 19226 636
rect 19238 602 19271 636
rect 19271 602 19290 636
rect 19302 602 19305 636
rect 19305 602 19343 636
rect 19343 602 19354 636
rect 19366 602 19377 636
rect 19377 602 19415 636
rect 19415 602 19418 636
rect 19430 602 19449 636
rect 19449 602 19482 636
rect 19494 602 19521 636
rect 19521 602 19546 636
rect 19174 593 19226 602
rect 19238 593 19290 602
rect 19302 593 19354 602
rect 19366 593 19418 602
rect 19430 593 19482 602
rect 19494 593 19546 602
rect 19558 636 19610 645
rect 19558 602 19559 636
rect 19559 602 19593 636
rect 19593 602 19610 636
rect 19558 593 19610 602
rect 19622 636 19674 645
rect 19622 602 19631 636
rect 19631 602 19665 636
rect 19665 602 19674 636
rect 19622 593 19674 602
rect 19686 636 19738 645
rect 19686 602 19703 636
rect 19703 602 19737 636
rect 19737 602 19738 636
rect 19686 593 19738 602
rect 19750 636 19802 645
rect 19814 636 19866 645
rect 19878 636 19930 645
rect 19942 636 19994 645
rect 20006 636 20058 645
rect 20070 636 20122 645
rect 19750 602 19775 636
rect 19775 602 19802 636
rect 19814 602 19847 636
rect 19847 602 19866 636
rect 19878 602 19881 636
rect 19881 602 19919 636
rect 19919 602 19930 636
rect 19942 602 19953 636
rect 19953 602 19991 636
rect 19991 602 19994 636
rect 20006 602 20025 636
rect 20025 602 20058 636
rect 20070 602 20097 636
rect 20097 602 20122 636
rect 19750 593 19802 602
rect 19814 593 19866 602
rect 19878 593 19930 602
rect 19942 593 19994 602
rect 20006 593 20058 602
rect 20070 593 20122 602
rect 20134 636 20186 645
rect 20134 602 20135 636
rect 20135 602 20169 636
rect 20169 602 20186 636
rect 20134 593 20186 602
rect 20198 636 20250 645
rect 20198 602 20207 636
rect 20207 602 20241 636
rect 20241 602 20250 636
rect 20198 593 20250 602
rect 20262 636 20314 645
rect 20262 602 20279 636
rect 20279 602 20313 636
rect 20313 602 20314 636
rect 20262 593 20314 602
rect 20326 636 20378 645
rect 20390 636 20442 645
rect 20454 636 20506 645
rect 20518 636 20570 645
rect 20582 636 20634 645
rect 20646 636 20698 645
rect 20326 602 20351 636
rect 20351 602 20378 636
rect 20390 602 20423 636
rect 20423 602 20442 636
rect 20454 602 20457 636
rect 20457 602 20495 636
rect 20495 602 20506 636
rect 20518 602 20529 636
rect 20529 602 20567 636
rect 20567 602 20570 636
rect 20582 602 20601 636
rect 20601 602 20634 636
rect 20646 602 20673 636
rect 20673 602 20698 636
rect 20326 593 20378 602
rect 20390 593 20442 602
rect 20454 593 20506 602
rect 20518 593 20570 602
rect 20582 593 20634 602
rect 20646 593 20698 602
rect 20710 636 20762 645
rect 20710 602 20711 636
rect 20711 602 20745 636
rect 20745 602 20762 636
rect 20710 593 20762 602
rect 20774 636 20826 645
rect 20774 602 20783 636
rect 20783 602 20817 636
rect 20817 602 20826 636
rect 20774 593 20826 602
rect 20838 636 20890 645
rect 20838 602 20855 636
rect 20855 602 20889 636
rect 20889 602 20890 636
rect 20838 593 20890 602
rect 20902 636 20954 645
rect 20966 636 21018 645
rect 21030 636 21082 645
rect 21094 636 21146 645
rect 21158 636 21210 645
rect 21222 636 21274 645
rect 20902 602 20927 636
rect 20927 602 20954 636
rect 20966 602 20999 636
rect 20999 602 21018 636
rect 21030 602 21033 636
rect 21033 602 21071 636
rect 21071 602 21082 636
rect 21094 602 21105 636
rect 21105 602 21143 636
rect 21143 602 21146 636
rect 21158 602 21177 636
rect 21177 602 21210 636
rect 21222 602 21249 636
rect 21249 602 21274 636
rect 20902 593 20954 602
rect 20966 593 21018 602
rect 21030 593 21082 602
rect 21094 593 21146 602
rect 21158 593 21210 602
rect 21222 593 21274 602
rect 21286 636 21338 645
rect 21286 602 21287 636
rect 21287 602 21321 636
rect 21321 602 21338 636
rect 21286 593 21338 602
rect 21350 636 21402 645
rect 21350 602 21359 636
rect 21359 602 21393 636
rect 21393 602 21402 636
rect 21350 593 21402 602
rect 21414 636 21466 645
rect 21414 602 21431 636
rect 21431 602 21465 636
rect 21465 602 21466 636
rect 21414 593 21466 602
rect 21478 636 21530 645
rect 21542 636 21594 645
rect 21606 636 21658 645
rect 21670 636 21722 645
rect 21734 636 21786 645
rect 21798 636 21850 645
rect 21478 602 21503 636
rect 21503 602 21530 636
rect 21542 602 21575 636
rect 21575 602 21594 636
rect 21606 602 21609 636
rect 21609 602 21647 636
rect 21647 602 21658 636
rect 21670 602 21681 636
rect 21681 602 21719 636
rect 21719 602 21722 636
rect 21734 602 21753 636
rect 21753 602 21786 636
rect 21798 602 21825 636
rect 21825 602 21850 636
rect 21478 593 21530 602
rect 21542 593 21594 602
rect 21606 593 21658 602
rect 21670 593 21722 602
rect 21734 593 21786 602
rect 21798 593 21850 602
rect 21862 636 21914 645
rect 21862 602 21863 636
rect 21863 602 21897 636
rect 21897 602 21914 636
rect 21862 593 21914 602
rect 21926 636 21978 645
rect 21926 602 21935 636
rect 21935 602 21969 636
rect 21969 602 21978 636
rect 21926 593 21978 602
rect 20694 473 20746 525
rect 20760 473 20812 525
rect 20826 473 20878 525
rect 20892 473 20944 525
rect 20957 473 21009 525
rect 21022 473 21074 525
rect 20694 409 20746 461
rect 20760 409 20812 461
rect 20826 409 20878 461
rect 20892 409 20944 461
rect 20957 409 21009 461
rect 21022 409 21074 461
rect 20694 345 20746 397
rect 20760 345 20812 397
rect 20826 345 20878 397
rect 20892 345 20944 397
rect 20957 345 21009 397
rect 21022 345 21074 397
rect 23407 473 23459 525
rect 23478 473 23530 525
rect 23549 473 23601 525
rect 23620 473 23672 525
rect 23691 473 23743 525
rect 23761 473 23813 525
rect 23831 473 23883 525
rect 23901 473 23953 525
rect 23971 473 24023 525
rect 24041 473 24093 525
rect 23407 409 23459 461
rect 23478 409 23530 461
rect 23549 409 23601 461
rect 23620 409 23672 461
rect 23691 409 23743 461
rect 23761 409 23813 461
rect 23831 409 23883 461
rect 23901 409 23953 461
rect 23971 409 24023 461
rect 24041 409 24093 461
rect 23407 345 23459 397
rect 23478 345 23530 397
rect 23549 345 23601 397
rect 23620 345 23672 397
rect 23691 345 23743 397
rect 23761 345 23813 397
rect 23831 345 23883 397
rect 23901 345 23953 397
rect 23971 345 24023 397
rect 24041 345 24093 397
<< metal2 >>
tri 22295 3032 22430 3167 se
rect 22430 3032 23308 3361
rect 19376 3028 23308 3032
rect 18581 2972 18590 3028
rect 18646 2972 18672 3028
rect 18728 2972 18754 3028
rect 18810 2972 18836 3028
rect 18892 2972 18918 3028
rect 18974 2972 19000 3028
rect 19056 2972 19082 3028
rect 19138 2972 19164 3028
rect 19220 2972 19247 3028
rect 19303 2972 19330 3028
rect 19386 2972 19413 3028
rect 19469 2972 23308 3028
rect 18581 2894 23308 2972
rect 18581 2838 18590 2894
rect 18646 2838 18672 2894
rect 18728 2838 18754 2894
rect 18810 2838 18836 2894
rect 18892 2838 18918 2894
rect 18974 2838 19000 2894
rect 19056 2838 19082 2894
rect 19138 2838 19164 2894
rect 19220 2838 19247 2894
rect 19303 2838 19330 2894
rect 19386 2838 19413 2894
rect 19469 2838 23308 2894
rect 19376 2834 23308 2838
tri 22330 2734 22430 2834 ne
rect 22430 2115 23308 2834
rect 22430 2063 22436 2115
rect 22488 2063 22504 2115
rect 22556 2063 22572 2115
rect 22624 2063 22640 2115
rect 22692 2063 22708 2115
rect 22760 2063 22776 2115
rect 22828 2063 22844 2115
rect 22896 2063 22912 2115
rect 22964 2063 22980 2115
rect 23032 2063 23048 2115
rect 23100 2063 23116 2115
rect 23168 2063 23183 2115
rect 23235 2063 23250 2115
rect 23302 2063 23308 2115
rect 22236 2055 22288 2061
rect 22236 1991 22288 2003
rect 22236 1927 22288 1939
rect 22236 1863 22288 1875
rect 22236 1799 22288 1811
rect 22236 1735 22288 1747
rect 22236 1671 22288 1683
rect 22236 1607 22288 1619
rect 22236 1543 22288 1555
rect 22236 1479 22288 1491
rect 22236 1415 22288 1427
rect 22236 1351 22288 1363
rect 22236 1287 22288 1299
rect 7714 1269 7723 1271
rect 7779 1269 7806 1271
rect 7862 1269 7888 1271
rect 7944 1269 7970 1271
rect 8026 1269 8052 1271
rect 8108 1269 8117 1271
rect 8645 1269 8654 1271
rect 8710 1269 8737 1271
rect 8793 1269 8819 1271
rect 8875 1269 8901 1271
rect 8957 1269 8983 1271
rect 9039 1269 9048 1271
rect 14202 1270 14211 1271
rect 14267 1270 14294 1271
rect 14350 1270 14376 1271
rect 14432 1270 14458 1271
rect 14514 1270 14540 1271
rect 14596 1270 14605 1271
rect 15129 1270 15138 1271
rect 15194 1270 15221 1271
rect 15277 1270 15303 1271
rect 15359 1270 15385 1271
rect 15441 1270 15467 1271
rect 15523 1270 15532 1271
rect 20767 1270 20776 1271
rect 20832 1270 20859 1271
rect 20915 1270 20942 1271
rect 20998 1270 21024 1271
rect 21080 1270 21089 1271
rect 7610 1217 7616 1269
rect 7668 1217 7681 1269
rect 7798 1217 7806 1269
rect 7863 1217 7876 1269
rect 8123 1217 8136 1269
rect 8188 1217 8201 1269
rect 8253 1217 8266 1269
rect 8318 1217 8331 1269
rect 8383 1217 8396 1269
rect 8448 1217 8461 1269
rect 8513 1217 8526 1269
rect 8578 1217 8591 1269
rect 8643 1217 8654 1269
rect 8710 1217 8721 1269
rect 8968 1217 8981 1269
rect 9039 1217 9046 1269
rect 9098 1217 9111 1269
rect 9163 1217 9176 1269
rect 9228 1217 9241 1269
rect 9293 1217 9306 1269
rect 9358 1217 9371 1269
rect 9423 1217 9436 1269
rect 9488 1217 9501 1269
rect 9553 1217 9566 1269
rect 9618 1217 9631 1269
rect 9683 1217 9696 1269
rect 9748 1217 9761 1269
rect 9813 1217 9826 1269
rect 9878 1217 9891 1269
rect 9943 1217 9956 1269
rect 10008 1217 10021 1269
rect 10073 1217 10086 1269
rect 10138 1217 10151 1269
rect 10203 1217 10216 1269
rect 10268 1217 10281 1269
rect 10333 1217 10346 1269
rect 10398 1217 10411 1269
rect 10463 1217 10476 1269
rect 10528 1217 10541 1269
rect 10593 1217 10606 1269
rect 10658 1217 10671 1269
rect 10723 1217 10736 1269
rect 10788 1217 10800 1269
rect 10852 1217 10864 1269
rect 10916 1217 10928 1269
rect 10980 1217 10992 1269
rect 11044 1217 11056 1269
rect 11108 1217 11120 1269
rect 11172 1217 11184 1269
rect 11236 1217 11248 1269
rect 11300 1217 11312 1269
rect 11364 1217 11376 1269
rect 11428 1217 11440 1269
rect 11492 1217 11504 1269
rect 11556 1217 11568 1269
rect 11620 1217 11632 1269
rect 11684 1217 11696 1269
rect 11748 1217 11760 1269
rect 11812 1217 11824 1269
rect 11876 1217 11882 1269
rect 12588 1218 12594 1270
rect 12646 1218 12659 1270
rect 12711 1218 12724 1270
rect 12776 1218 12789 1270
rect 12841 1218 12854 1270
rect 12906 1218 12919 1270
rect 12971 1218 12984 1270
rect 13036 1218 13049 1270
rect 13101 1218 13114 1270
rect 13166 1218 13179 1270
rect 13231 1218 13244 1270
rect 13296 1218 13309 1270
rect 13361 1218 13374 1270
rect 13426 1218 13439 1270
rect 13491 1218 13504 1270
rect 13556 1218 13569 1270
rect 13621 1218 13633 1270
rect 13685 1218 13697 1270
rect 13749 1218 13761 1270
rect 13813 1218 13825 1270
rect 13877 1218 13889 1270
rect 13941 1218 13953 1270
rect 14005 1218 14017 1270
rect 14069 1218 14081 1270
rect 14133 1218 14145 1270
rect 14197 1218 14209 1270
rect 14267 1218 14273 1270
rect 14453 1218 14458 1270
rect 14517 1218 14529 1270
rect 14645 1218 14657 1270
rect 14709 1218 14721 1270
rect 14773 1218 14785 1270
rect 14837 1218 14849 1270
rect 14901 1218 14913 1270
rect 14965 1218 14977 1270
rect 15029 1218 15041 1270
rect 15093 1218 15105 1270
rect 15285 1218 15297 1270
rect 15359 1218 15361 1270
rect 15541 1218 15553 1270
rect 15605 1218 15617 1270
rect 15669 1218 15681 1270
rect 15733 1218 15745 1270
rect 15797 1218 15809 1270
rect 15861 1218 15873 1270
rect 15925 1218 15937 1270
rect 15989 1218 16001 1270
rect 16053 1218 16065 1270
rect 16117 1218 16129 1270
rect 16181 1218 16193 1270
rect 16245 1218 16257 1270
rect 16309 1218 16321 1270
rect 16373 1218 16385 1270
rect 16437 1218 16449 1270
rect 16501 1218 16513 1270
rect 16565 1218 16577 1270
rect 16629 1218 16641 1270
rect 16693 1218 16705 1270
rect 16757 1218 16769 1270
rect 16821 1218 16833 1270
rect 16885 1218 16897 1270
rect 16949 1218 16961 1270
rect 17013 1218 17025 1270
rect 17077 1218 17089 1270
rect 17141 1218 17153 1270
rect 17205 1218 17217 1270
rect 17269 1218 17281 1270
rect 17333 1218 17345 1270
rect 17397 1218 17409 1270
rect 17461 1218 17473 1270
rect 17525 1218 17537 1270
rect 17589 1218 17601 1270
rect 17653 1218 17665 1270
rect 17717 1218 17729 1270
rect 17781 1218 17793 1270
rect 17845 1218 17857 1270
rect 17909 1218 17921 1270
rect 17973 1218 17985 1270
rect 18037 1218 18049 1270
rect 18101 1218 18113 1270
rect 18165 1218 18177 1270
rect 18229 1218 18241 1270
rect 18293 1218 18305 1270
rect 18357 1218 18369 1270
rect 18421 1218 18433 1270
rect 18485 1218 18497 1270
rect 18549 1218 18561 1270
rect 18613 1218 18625 1270
rect 18677 1218 18689 1270
rect 18741 1218 18753 1270
rect 18805 1218 18817 1270
rect 18869 1218 18881 1270
rect 18933 1218 18945 1270
rect 18997 1218 19009 1270
rect 19061 1218 19073 1270
rect 19125 1218 19137 1270
rect 19189 1218 19201 1270
rect 19253 1218 19265 1270
rect 19317 1218 19329 1270
rect 19381 1218 19393 1270
rect 19445 1218 19457 1270
rect 19509 1218 19521 1270
rect 19573 1218 19585 1270
rect 19637 1218 19649 1270
rect 19701 1218 19713 1270
rect 19765 1218 19777 1270
rect 19829 1218 19841 1270
rect 19893 1218 19905 1270
rect 19957 1218 19969 1270
rect 20021 1218 20033 1270
rect 20085 1218 20097 1270
rect 20149 1218 20161 1270
rect 20213 1218 20225 1270
rect 20277 1218 20289 1270
rect 20341 1218 20353 1270
rect 20405 1218 20417 1270
rect 20469 1218 20481 1270
rect 20533 1218 20545 1270
rect 20597 1218 20609 1270
rect 20661 1218 20673 1270
rect 20725 1218 20737 1270
rect 20853 1218 20859 1270
rect 20917 1218 20929 1270
rect 21109 1218 21121 1270
rect 21173 1218 21185 1270
rect 21237 1218 21249 1270
rect 21301 1218 21313 1270
rect 21365 1218 21377 1270
rect 21429 1218 21441 1270
rect 21493 1218 21505 1270
rect 21557 1218 21569 1270
rect 21621 1218 21633 1270
rect 21685 1218 21697 1270
rect 21749 1218 21761 1270
rect 21813 1218 21825 1270
rect 21877 1218 21889 1270
rect 21941 1218 21947 1270
rect 22236 1223 22288 1235
rect 7714 1215 7723 1217
rect 7779 1215 7806 1217
rect 7862 1215 7888 1217
rect 7944 1215 7970 1217
rect 8026 1215 8052 1217
rect 8108 1215 8117 1217
rect 8645 1215 8654 1217
rect 8710 1215 8737 1217
rect 8793 1215 8819 1217
rect 8875 1215 8901 1217
rect 8957 1215 8983 1217
rect 9039 1215 9048 1217
rect 14202 1215 14211 1218
rect 14267 1215 14294 1218
rect 14350 1215 14376 1218
rect 14432 1215 14458 1218
rect 14514 1215 14540 1218
rect 14596 1215 14605 1218
rect 15129 1215 15138 1218
rect 15194 1215 15221 1218
rect 15277 1215 15303 1218
rect 15359 1215 15385 1218
rect 15441 1215 15467 1218
rect 15523 1215 15532 1218
rect 20767 1215 20776 1218
rect 20832 1215 20859 1218
rect 20915 1215 20942 1218
rect 20998 1215 21024 1218
rect 21080 1215 21089 1218
rect 22236 1159 22288 1171
tri 10258 1113 10260 1115 se
rect 10260 1113 10269 1115
rect 10325 1113 10351 1115
rect 10407 1113 10433 1115
rect 10489 1113 10515 1115
rect 10571 1113 10597 1115
rect 10653 1113 10679 1115
rect 10735 1113 10760 1115
rect 10816 1113 10841 1115
rect 10897 1113 10922 1115
rect 10978 1113 11003 1115
rect 11059 1113 11084 1115
rect 11140 1113 11149 1115
tri 11149 1113 11151 1115 sw
tri 12099 1113 12101 1115 se
rect 12101 1113 12110 1115
rect 12166 1113 12192 1115
rect 12248 1113 12274 1115
rect 12330 1113 12356 1115
rect 12412 1113 12438 1115
rect 12494 1113 12520 1115
rect 12576 1113 12601 1115
rect 12657 1113 12682 1115
rect 12738 1113 12763 1115
rect 12819 1113 12844 1115
rect 12900 1113 12925 1115
rect 12981 1113 12990 1115
tri 12990 1113 12992 1115 sw
tri 16742 1113 16744 1115 se
rect 16744 1113 16753 1115
rect 16809 1113 16835 1115
rect 16891 1113 16917 1115
rect 16973 1113 16999 1115
rect 17055 1113 17081 1115
rect 17137 1113 17163 1115
rect 17219 1113 17244 1115
rect 17300 1113 17325 1115
rect 17381 1113 17406 1115
rect 17462 1113 17487 1115
rect 17543 1113 17568 1115
rect 17624 1113 17633 1115
tri 17633 1113 17635 1115 sw
tri 18583 1113 18585 1115 se
rect 18585 1113 18594 1115
rect 18650 1113 18676 1115
rect 18732 1113 18758 1115
rect 18814 1113 18840 1115
rect 18896 1113 18922 1115
rect 18978 1113 19004 1115
rect 19060 1113 19085 1115
rect 19141 1113 19166 1115
rect 19222 1113 19247 1115
rect 19303 1113 19328 1115
rect 19384 1113 19409 1115
rect 19465 1113 19474 1115
tri 19474 1113 19476 1115 sw
rect 7610 1061 7616 1113
rect 7668 1061 7681 1113
rect 7733 1061 7746 1113
rect 7798 1061 7811 1113
rect 7863 1061 7876 1113
rect 7928 1061 7941 1113
rect 7993 1061 8006 1113
rect 8058 1061 8071 1113
rect 8123 1061 8136 1113
rect 8188 1061 8201 1113
rect 8253 1061 8266 1113
rect 8318 1061 8331 1113
rect 8383 1061 8396 1113
rect 8448 1061 8461 1113
rect 8513 1061 8526 1113
rect 8578 1061 8591 1113
rect 8643 1061 8656 1113
rect 8708 1061 8721 1113
rect 8773 1061 8786 1113
rect 8838 1061 8851 1113
rect 8903 1061 8916 1113
rect 8968 1061 8981 1113
rect 9033 1061 9046 1113
rect 9098 1061 9111 1113
rect 9163 1061 9176 1113
rect 9228 1061 9241 1113
rect 9293 1061 9306 1113
rect 9358 1061 9371 1113
rect 9423 1061 9436 1113
rect 9488 1061 9501 1113
rect 9553 1061 9566 1113
rect 9618 1061 9631 1113
rect 9683 1061 9696 1113
rect 9748 1061 9761 1113
rect 9813 1061 9826 1113
rect 9878 1061 9891 1113
rect 9943 1061 9956 1113
rect 10008 1061 10021 1113
rect 10073 1061 10086 1113
rect 10138 1061 10151 1113
rect 10203 1061 10216 1113
rect 10268 1061 10269 1113
rect 10333 1061 10346 1113
rect 10407 1061 10411 1113
rect 10593 1061 10597 1113
rect 10658 1061 10671 1113
rect 10735 1061 10736 1113
rect 10916 1061 10922 1113
rect 10980 1061 10992 1113
rect 11172 1061 11184 1113
rect 11236 1061 11248 1113
rect 11300 1061 11312 1113
rect 11364 1061 11376 1113
rect 11428 1061 11440 1113
rect 11492 1061 11504 1113
rect 11556 1061 11568 1113
rect 11620 1061 11632 1113
rect 11684 1061 11696 1113
rect 11748 1061 11760 1113
rect 11812 1061 11824 1113
rect 11876 1061 11882 1113
rect 12016 1061 12022 1113
rect 12074 1061 12087 1113
rect 12269 1061 12274 1113
rect 12334 1061 12347 1113
rect 12594 1061 12601 1113
rect 12659 1061 12672 1113
rect 12917 1061 12925 1113
rect 12981 1061 12993 1113
rect 13045 1061 13057 1113
rect 13109 1061 13121 1113
rect 13173 1061 13185 1113
rect 13237 1061 13249 1113
rect 13301 1061 13313 1113
rect 13365 1061 13377 1113
rect 13429 1061 13441 1113
rect 13493 1061 13505 1113
rect 13557 1061 13569 1113
rect 13621 1061 13633 1113
rect 13685 1061 13697 1113
rect 13749 1061 13761 1113
rect 13813 1061 13825 1113
rect 13877 1061 13889 1113
rect 13941 1061 13953 1113
rect 14005 1061 14017 1113
rect 14069 1061 14081 1113
rect 14133 1061 14145 1113
rect 14197 1061 14209 1113
rect 14261 1061 14273 1113
rect 14325 1061 14337 1113
rect 14389 1061 14401 1113
rect 14453 1061 14465 1113
rect 14517 1061 14529 1113
rect 14581 1061 14593 1113
rect 14645 1061 14657 1113
rect 14709 1061 14721 1113
rect 14773 1061 14785 1113
rect 14837 1061 14849 1113
rect 14901 1061 14913 1113
rect 14965 1061 14977 1113
rect 15029 1061 15041 1113
rect 15093 1061 15105 1113
rect 15157 1061 15169 1113
rect 15221 1061 15233 1113
rect 15285 1061 15297 1113
rect 15349 1061 15361 1113
rect 15413 1061 15425 1113
rect 15477 1061 15489 1113
rect 15541 1061 15553 1113
rect 15605 1061 15617 1113
rect 15669 1061 15681 1113
rect 15733 1061 15745 1113
rect 15797 1061 15809 1113
rect 15861 1061 15873 1113
rect 15925 1061 15937 1113
rect 15989 1061 16001 1113
rect 16053 1061 16065 1113
rect 16117 1061 16129 1113
rect 16181 1061 16193 1113
rect 16245 1061 16257 1113
rect 16309 1061 16321 1113
rect 16373 1061 16385 1113
rect 16437 1061 16449 1113
rect 16501 1061 16513 1113
rect 16565 1061 16577 1113
rect 16629 1061 16641 1113
rect 16693 1061 16705 1113
rect 16821 1061 16833 1113
rect 16891 1061 16897 1113
rect 17077 1061 17081 1113
rect 17141 1061 17153 1113
rect 17397 1061 17406 1113
rect 17462 1061 17473 1113
rect 17653 1061 17665 1113
rect 17717 1061 17729 1113
rect 17781 1061 17793 1113
rect 17845 1061 17857 1113
rect 17909 1061 17921 1113
rect 17973 1061 17985 1113
rect 18037 1061 18049 1113
rect 18101 1061 18113 1113
rect 18165 1061 18177 1113
rect 18229 1061 18241 1113
rect 18293 1061 18305 1113
rect 18357 1061 18369 1113
rect 18421 1061 18433 1113
rect 18485 1061 18497 1113
rect 18549 1061 18561 1113
rect 18741 1061 18753 1113
rect 18814 1061 18817 1113
rect 18997 1061 19004 1113
rect 19061 1061 19073 1113
rect 19317 1061 19328 1113
rect 19384 1061 19393 1113
rect 19509 1061 19521 1113
rect 19573 1061 19585 1113
rect 19637 1061 19649 1113
rect 19701 1061 19713 1113
rect 19765 1061 19777 1113
rect 19829 1061 19841 1113
rect 19893 1061 19905 1113
rect 19957 1061 19969 1113
rect 20021 1061 20033 1113
rect 20085 1061 20097 1113
rect 20149 1061 20161 1113
rect 20213 1061 20225 1113
rect 20277 1061 20289 1113
rect 20341 1061 20353 1113
rect 20405 1061 20417 1113
rect 20469 1061 20481 1113
rect 20533 1061 20545 1113
rect 20597 1061 20609 1113
rect 20661 1061 20673 1113
rect 20725 1061 20737 1113
rect 20789 1061 20801 1113
rect 20853 1061 20865 1113
rect 20917 1061 20929 1113
rect 20981 1061 20993 1113
rect 21045 1061 21057 1113
rect 21109 1061 21121 1113
rect 21173 1061 21185 1113
rect 21237 1061 21249 1113
rect 21301 1061 21313 1113
rect 21365 1061 21377 1113
rect 21429 1061 21441 1113
rect 21493 1061 21505 1113
rect 21557 1061 21569 1113
rect 21621 1061 21633 1113
rect 21685 1061 21697 1113
rect 21749 1061 21761 1113
rect 21813 1061 21825 1113
rect 21877 1061 21889 1113
rect 21941 1061 21947 1113
rect 22236 1095 22288 1107
tri 10258 1059 10260 1061 ne
rect 10260 1059 10269 1061
rect 10325 1059 10351 1061
rect 10407 1059 10433 1061
rect 10489 1059 10515 1061
rect 10571 1059 10597 1061
rect 10653 1059 10679 1061
rect 10735 1059 10760 1061
rect 10816 1059 10841 1061
rect 10897 1059 10922 1061
rect 10978 1059 11003 1061
rect 11059 1059 11084 1061
rect 11140 1059 11149 1061
tri 11149 1059 11151 1061 nw
tri 12099 1059 12101 1061 ne
rect 12101 1059 12110 1061
rect 12166 1059 12192 1061
rect 12248 1059 12274 1061
rect 12330 1059 12356 1061
rect 12412 1059 12438 1061
rect 12494 1059 12520 1061
rect 12576 1059 12601 1061
rect 12657 1059 12682 1061
rect 12738 1059 12763 1061
rect 12819 1059 12844 1061
rect 12900 1059 12925 1061
rect 12981 1059 12990 1061
tri 12990 1059 12992 1061 nw
tri 16742 1059 16744 1061 ne
rect 16744 1059 16753 1061
rect 16809 1059 16835 1061
rect 16891 1059 16917 1061
rect 16973 1059 16999 1061
rect 17055 1059 17081 1061
rect 17137 1059 17163 1061
rect 17219 1059 17244 1061
rect 17300 1059 17325 1061
rect 17381 1059 17406 1061
rect 17462 1059 17487 1061
rect 17543 1059 17568 1061
rect 17624 1059 17633 1061
tri 17633 1059 17635 1061 nw
tri 18583 1059 18585 1061 ne
rect 18585 1059 18594 1061
rect 18650 1059 18676 1061
rect 18732 1059 18758 1061
rect 18814 1059 18840 1061
rect 18896 1059 18922 1061
rect 18978 1059 19004 1061
rect 19060 1059 19085 1061
rect 19141 1059 19166 1061
rect 19222 1059 19247 1061
rect 19303 1059 19328 1061
rect 19384 1059 19409 1061
rect 19465 1059 19474 1061
tri 19474 1059 19476 1061 nw
rect 22236 1031 22288 1043
rect 22236 967 22288 979
rect 7714 957 7723 959
rect 7779 957 7806 959
rect 7862 957 7888 959
rect 7944 957 7970 959
rect 8026 957 8052 959
rect 8108 957 8117 959
rect 8645 957 8654 959
rect 8710 957 8737 959
rect 8793 957 8819 959
rect 8875 957 8901 959
rect 8957 957 8983 959
rect 9039 957 9048 959
rect 14198 957 14207 959
rect 14263 957 14290 959
rect 14346 957 14372 959
rect 14428 957 14454 959
rect 14510 957 14536 959
rect 14592 957 14601 959
rect 15129 957 15138 959
rect 15194 957 15221 959
rect 15277 957 15303 959
rect 15359 957 15385 959
rect 15441 957 15467 959
rect 15523 957 15532 959
rect 20767 957 20776 959
rect 20832 957 20858 959
rect 20914 957 20939 959
rect 20995 957 21020 959
rect 21076 957 21085 959
rect 7610 905 7616 957
rect 7668 905 7681 957
rect 7798 905 7806 957
rect 7863 905 7876 957
rect 8123 905 8136 957
rect 8188 905 8201 957
rect 8253 905 8266 957
rect 8318 905 8331 957
rect 8383 905 8396 957
rect 8448 905 8461 957
rect 8513 905 8526 957
rect 8578 905 8591 957
rect 8643 905 8654 957
rect 8710 905 8721 957
rect 8968 905 8981 957
rect 9039 905 9046 957
rect 9098 905 9111 957
rect 9163 905 9176 957
rect 9228 905 9241 957
rect 9293 905 9306 957
rect 9358 905 9371 957
rect 9423 905 9436 957
rect 9488 905 9501 957
rect 9553 905 9566 957
rect 9618 905 9631 957
rect 9683 905 9696 957
rect 9748 905 9761 957
rect 9813 905 9826 957
rect 9878 905 9891 957
rect 9943 905 9956 957
rect 10008 905 10021 957
rect 10073 905 10086 957
rect 10138 905 10151 957
rect 10203 905 10216 957
rect 10268 905 10281 957
rect 10333 905 10346 957
rect 10398 905 10411 957
rect 10463 905 10476 957
rect 10528 905 10541 957
rect 10593 905 10606 957
rect 10658 905 10671 957
rect 10723 905 10736 957
rect 10788 905 10800 957
rect 10852 905 10864 957
rect 10916 905 10928 957
rect 10980 905 10992 957
rect 11044 905 11056 957
rect 11108 905 11120 957
rect 11172 905 11184 957
rect 11236 905 11248 957
rect 11300 905 11312 957
rect 11364 905 11376 957
rect 11428 905 11440 957
rect 11492 905 11504 957
rect 11556 905 11568 957
rect 11620 905 11632 957
rect 11684 905 11696 957
rect 11748 905 11760 957
rect 11812 905 11824 957
rect 11876 905 11882 957
rect 12016 905 12022 957
rect 12074 905 12087 957
rect 12139 905 12152 957
rect 12204 905 12217 957
rect 12269 905 12282 957
rect 12334 905 12347 957
rect 12399 905 12412 957
rect 12464 905 12477 957
rect 12529 905 12542 957
rect 12594 905 12607 957
rect 12659 905 12672 957
rect 12724 905 12737 957
rect 12789 905 12802 957
rect 12854 905 12867 957
rect 12919 905 12932 957
rect 12984 905 12997 957
rect 13049 905 13062 957
rect 13114 905 13127 957
rect 13179 905 13192 957
rect 13244 905 13257 957
rect 13309 905 13322 957
rect 13374 905 13387 957
rect 13439 905 13452 957
rect 13504 905 13517 957
rect 13569 905 13582 957
rect 13634 905 13647 957
rect 13699 905 13712 957
rect 13764 905 13777 957
rect 13829 905 13842 957
rect 13894 905 13907 957
rect 13959 905 13972 957
rect 14024 905 14037 957
rect 14089 905 14102 957
rect 14154 905 14167 957
rect 14284 905 14290 957
rect 14349 905 14362 957
rect 14609 905 14622 957
rect 14674 905 14686 957
rect 14738 905 14750 957
rect 14802 905 14814 957
rect 14866 905 14878 957
rect 14930 905 14942 957
rect 14994 905 15006 957
rect 15058 905 15070 957
rect 15122 905 15134 957
rect 15194 905 15198 957
rect 15378 905 15385 957
rect 15442 905 15454 957
rect 15570 905 15582 957
rect 15634 905 15646 957
rect 15698 905 15710 957
rect 15762 905 15774 957
rect 15826 905 15838 957
rect 15890 905 15902 957
rect 15954 905 15966 957
rect 16018 905 16030 957
rect 16082 905 16094 957
rect 16146 905 16158 957
rect 16210 905 16222 957
rect 16274 905 16286 957
rect 16338 905 16350 957
rect 16402 905 16414 957
rect 16466 905 16478 957
rect 16530 905 16542 957
rect 16594 905 16606 957
rect 16658 905 16670 957
rect 16722 905 16734 957
rect 16786 905 16798 957
rect 16850 905 16862 957
rect 16914 905 16926 957
rect 16978 905 16990 957
rect 17042 905 17054 957
rect 17106 905 17118 957
rect 17170 905 17182 957
rect 17234 905 17246 957
rect 17298 905 17310 957
rect 17362 905 17374 957
rect 17426 905 17438 957
rect 17490 905 17502 957
rect 17554 905 17566 957
rect 17618 905 17630 957
rect 17682 905 17694 957
rect 17746 905 17758 957
rect 17810 905 17822 957
rect 17874 905 17886 957
rect 17938 905 17950 957
rect 18002 905 18014 957
rect 18066 905 18078 957
rect 18130 905 18142 957
rect 18194 905 18206 957
rect 18258 905 18270 957
rect 18322 905 18334 957
rect 18386 905 18398 957
rect 18450 905 18462 957
rect 18514 905 18526 957
rect 18578 905 18590 957
rect 18642 905 18654 957
rect 18706 905 18718 957
rect 18770 905 18782 957
rect 18834 905 18846 957
rect 18898 905 18910 957
rect 18962 905 18974 957
rect 19026 905 19038 957
rect 19090 905 19102 957
rect 19154 905 19166 957
rect 19218 905 19230 957
rect 19282 905 19294 957
rect 19346 905 19358 957
rect 19410 905 19422 957
rect 19474 905 19486 957
rect 19538 905 19550 957
rect 19602 905 19614 957
rect 19666 905 19678 957
rect 19730 905 19742 957
rect 19794 905 19806 957
rect 19858 905 19870 957
rect 19922 905 19934 957
rect 19986 905 19998 957
rect 20050 905 20062 957
rect 20114 905 20126 957
rect 20178 905 20190 957
rect 20242 905 20254 957
rect 20306 905 20318 957
rect 20370 905 20382 957
rect 20434 905 20446 957
rect 20498 905 20510 957
rect 20562 905 20574 957
rect 20626 905 20638 957
rect 20690 905 20702 957
rect 20754 905 20766 957
rect 21010 905 21020 957
rect 21076 905 21086 957
rect 21138 905 21150 957
rect 21202 905 21214 957
rect 21266 905 21278 957
rect 21330 905 21342 957
rect 21394 905 21406 957
rect 21458 905 21470 957
rect 21522 905 21534 957
rect 21586 905 21598 957
rect 21650 905 21662 957
rect 21714 905 21726 957
rect 21778 905 21790 957
rect 21842 905 21854 957
rect 21906 905 21918 957
rect 21970 905 21976 957
rect 7714 903 7723 905
rect 7779 903 7806 905
rect 7862 903 7888 905
rect 7944 903 7970 905
rect 8026 903 8052 905
rect 8108 903 8117 905
rect 8645 903 8654 905
rect 8710 903 8737 905
rect 8793 903 8819 905
rect 8875 903 8901 905
rect 8957 903 8983 905
rect 9039 903 9048 905
rect 14198 903 14207 905
rect 14263 903 14290 905
rect 14346 903 14372 905
rect 14428 903 14454 905
rect 14510 903 14536 905
rect 14592 903 14601 905
rect 15129 903 15138 905
rect 15194 903 15221 905
rect 15277 903 15303 905
rect 15359 903 15385 905
rect 15441 903 15467 905
rect 15523 903 15532 905
rect 20767 903 20776 905
rect 20832 903 20858 905
rect 20914 903 20939 905
rect 20995 903 21020 905
rect 21076 903 21085 905
rect 22236 902 22288 915
rect 22236 837 22288 850
tri 5615 827 5617 829 se
rect 5617 827 5626 829
rect 5682 827 5714 829
rect 5770 827 5802 829
rect 5858 827 5890 829
rect 5946 827 5978 829
rect 6034 827 6066 829
rect 1539 775 1545 827
rect 1597 775 1610 827
rect 1662 775 1675 827
rect 1727 775 1740 827
rect 1792 775 1805 827
rect 1857 775 1870 827
rect 1922 775 1935 827
rect 1987 775 2000 827
rect 2052 775 2065 827
rect 2117 775 2130 827
rect 2182 775 2195 827
rect 2247 775 2260 827
rect 2312 775 2325 827
rect 2377 775 2390 827
rect 2442 775 2455 827
rect 2507 775 2520 827
rect 2572 775 2585 827
rect 2637 775 2650 827
rect 2702 775 2715 827
rect 2767 775 2780 827
rect 2832 775 2845 827
rect 2897 775 2910 827
rect 2962 775 2975 827
rect 3027 775 3040 827
rect 3092 775 3105 827
rect 3157 775 3170 827
rect 3222 775 3235 827
rect 3287 775 3300 827
rect 3352 775 3365 827
rect 3417 775 3430 827
rect 3482 775 3495 827
rect 3547 775 3560 827
rect 3612 775 3625 827
rect 3677 775 3690 827
rect 3742 775 3755 827
rect 3807 775 3820 827
rect 3872 775 3885 827
rect 3937 775 3950 827
rect 4002 775 4015 827
rect 4067 775 4080 827
rect 4132 775 4144 827
rect 4196 775 4208 827
rect 4260 775 4272 827
rect 4324 775 4336 827
rect 4388 775 4400 827
rect 4452 775 4464 827
rect 4516 775 4528 827
rect 4580 775 4592 827
rect 4644 775 4656 827
rect 4708 775 4720 827
rect 4772 775 4784 827
rect 4836 775 4848 827
rect 4900 775 4912 827
rect 4964 775 4976 827
rect 5028 775 5040 827
rect 5092 775 5104 827
rect 5156 775 5168 827
rect 5220 775 5232 827
rect 5284 775 5296 827
rect 5348 775 5360 827
rect 5412 775 5424 827
rect 5476 775 5488 827
rect 5540 775 5552 827
rect 5604 775 5616 827
rect 5796 775 5802 827
rect 5860 775 5872 827
rect 6052 775 6064 827
tri 5615 773 5617 775 ne
rect 5617 773 5626 775
rect 5682 773 5714 775
rect 5770 773 5802 775
rect 5858 773 5890 775
rect 5946 773 5978 775
rect 6034 773 6066 775
rect 6122 773 6153 829
rect 6209 773 6218 829
tri 10258 801 10260 803 se
rect 10260 801 10269 803
rect 10325 801 10351 803
rect 10407 801 10433 803
rect 10489 801 10515 803
rect 10571 801 10597 803
rect 10653 801 10679 803
rect 10735 801 10760 803
rect 10816 801 10841 803
rect 10897 801 10922 803
rect 10978 801 11003 803
rect 11059 801 11084 803
rect 11140 801 11149 803
tri 11149 801 11151 803 sw
tri 12099 801 12101 803 se
rect 12101 801 12110 803
rect 12166 801 12192 803
rect 12248 801 12274 803
rect 12330 801 12356 803
rect 12412 801 12438 803
rect 12494 801 12520 803
rect 12576 801 12601 803
rect 12657 801 12682 803
rect 12738 801 12763 803
rect 12819 801 12844 803
rect 12900 801 12925 803
rect 12981 801 12990 803
tri 12990 801 12992 803 sw
tri 16742 801 16744 803 se
rect 16744 801 16753 803
rect 16809 801 16835 803
rect 16891 801 16917 803
rect 16973 801 16999 803
rect 17055 801 17081 803
rect 17137 801 17163 803
rect 17219 801 17244 803
rect 17300 801 17325 803
rect 17381 801 17406 803
rect 17462 801 17487 803
rect 17543 801 17568 803
rect 17624 801 17633 803
tri 17633 801 17635 803 sw
tri 18583 801 18585 803 se
rect 18585 801 18594 803
rect 18650 801 18676 803
rect 18732 801 18758 803
rect 18814 801 18840 803
rect 18896 801 18922 803
rect 18978 801 19004 803
rect 19060 801 19085 803
rect 19141 801 19166 803
rect 19222 801 19247 803
rect 19303 801 19328 803
rect 19384 801 19409 803
rect 19465 801 19474 803
tri 19474 801 19476 803 sw
rect 7610 749 7616 801
rect 7668 749 7681 801
rect 7733 749 7746 801
rect 7798 749 7811 801
rect 7863 749 7876 801
rect 7928 749 7941 801
rect 7993 749 8006 801
rect 8058 749 8071 801
rect 8123 749 8136 801
rect 8188 749 8201 801
rect 8253 749 8266 801
rect 8318 749 8331 801
rect 8383 749 8396 801
rect 8448 749 8461 801
rect 8513 749 8526 801
rect 8578 749 8591 801
rect 8643 749 8656 801
rect 8708 749 8721 801
rect 8773 749 8786 801
rect 8838 749 8851 801
rect 8903 749 8916 801
rect 8968 749 8981 801
rect 9033 749 9046 801
rect 9098 749 9111 801
rect 9163 749 9176 801
rect 9228 749 9241 801
rect 9293 749 9306 801
rect 9358 749 9371 801
rect 9423 749 9436 801
rect 9488 749 9501 801
rect 9553 749 9566 801
rect 9618 749 9631 801
rect 9683 749 9696 801
rect 9748 749 9761 801
rect 9813 749 9826 801
rect 9878 749 9891 801
rect 9943 749 9956 801
rect 10008 749 10021 801
rect 10073 749 10086 801
rect 10138 749 10151 801
rect 10203 749 10216 801
rect 10268 749 10269 801
rect 10333 749 10346 801
rect 10407 749 10411 801
rect 10593 749 10597 801
rect 10658 749 10671 801
rect 10735 749 10736 801
rect 10916 749 10922 801
rect 10980 749 10992 801
rect 11172 749 11184 801
rect 11236 749 11248 801
rect 11300 749 11312 801
rect 11364 749 11376 801
rect 11428 749 11440 801
rect 11492 749 11504 801
rect 11556 749 11568 801
rect 11620 749 11632 801
rect 11684 749 11696 801
rect 11748 749 11760 801
rect 11812 749 11824 801
rect 11876 749 11882 801
rect 12016 749 12022 801
rect 12074 749 12087 801
rect 12269 749 12274 801
rect 12334 749 12347 801
rect 12594 749 12601 801
rect 12659 749 12672 801
rect 12919 749 12925 801
rect 12984 749 12997 801
rect 13049 749 13062 801
rect 13114 749 13127 801
rect 13179 749 13192 801
rect 13244 749 13257 801
rect 13309 749 13322 801
rect 13374 749 13387 801
rect 13439 749 13452 801
rect 13504 749 13517 801
rect 13569 749 13582 801
rect 13634 749 13647 801
rect 13699 749 13712 801
rect 13764 749 13777 801
rect 13829 749 13842 801
rect 13894 749 13907 801
rect 13959 749 13972 801
rect 14024 749 14037 801
rect 14089 749 14101 801
rect 14153 749 14165 801
rect 14217 749 14229 801
rect 14281 749 14293 801
rect 14345 749 14357 801
rect 14409 749 14421 801
rect 14473 749 14485 801
rect 14537 749 14549 801
rect 14601 749 14613 801
rect 14665 749 14677 801
rect 14729 749 14741 801
rect 14793 749 14805 801
rect 14857 749 14869 801
rect 14921 749 14933 801
rect 14985 749 14997 801
rect 15049 749 15061 801
rect 15113 749 15125 801
rect 15177 749 15189 801
rect 15241 749 15253 801
rect 15305 749 15317 801
rect 15369 749 15381 801
rect 15433 749 15445 801
rect 15497 749 15509 801
rect 15561 749 15573 801
rect 15625 749 15637 801
rect 15689 749 15701 801
rect 15753 749 15765 801
rect 15817 749 15829 801
rect 15881 749 15893 801
rect 15945 749 15957 801
rect 16009 749 16021 801
rect 16073 749 16085 801
rect 16137 749 16149 801
rect 16201 749 16213 801
rect 16265 749 16277 801
rect 16329 749 16341 801
rect 16393 749 16405 801
rect 16457 749 16469 801
rect 16521 749 16533 801
rect 16585 749 16597 801
rect 16649 749 16661 801
rect 16713 749 16725 801
rect 16905 749 16917 801
rect 16973 749 16981 801
rect 17161 749 17163 801
rect 17225 749 17237 801
rect 17300 749 17301 801
rect 17481 749 17487 801
rect 17545 749 17557 801
rect 17673 749 17685 801
rect 17737 749 17749 801
rect 17801 749 17813 801
rect 17865 749 17877 801
rect 17929 749 17941 801
rect 17993 749 18005 801
rect 18057 749 18069 801
rect 18121 749 18133 801
rect 18185 749 18197 801
rect 18249 749 18261 801
rect 18313 749 18325 801
rect 18377 749 18389 801
rect 18441 749 18453 801
rect 18505 749 18517 801
rect 18569 749 18581 801
rect 18825 749 18837 801
rect 18896 749 18901 801
rect 19081 749 19085 801
rect 19145 749 19157 801
rect 19401 749 19409 801
rect 19465 749 19477 801
rect 19529 749 19541 801
rect 19593 749 19605 801
rect 19657 749 19669 801
rect 19721 749 19733 801
rect 19785 749 19797 801
rect 19849 749 19861 801
rect 19913 749 19925 801
rect 19977 749 19989 801
rect 20041 749 20053 801
rect 20105 749 20117 801
rect 20169 749 20181 801
rect 20233 749 20245 801
rect 20297 749 20309 801
rect 20361 749 20373 801
rect 20425 749 20437 801
rect 20489 749 20501 801
rect 20553 749 20565 801
rect 20617 749 20629 801
rect 20681 749 20693 801
rect 20745 749 20757 801
rect 20809 749 20821 801
rect 20873 749 20885 801
rect 20937 749 20949 801
rect 21001 749 21013 801
rect 21065 749 21077 801
rect 21129 749 21141 801
rect 21193 749 21205 801
rect 21257 749 21269 801
rect 21321 749 21333 801
rect 21385 749 21397 801
rect 21449 749 21461 801
rect 21513 749 21525 801
rect 21577 749 21589 801
rect 21641 749 21653 801
rect 21705 749 21717 801
rect 21769 749 21781 801
rect 21833 749 21845 801
rect 21897 749 21909 801
rect 21961 749 21967 801
rect 22236 772 22288 785
tri 10258 747 10260 749 ne
rect 10260 747 10269 749
rect 10325 747 10351 749
rect 10407 747 10433 749
rect 10489 747 10515 749
rect 10571 747 10597 749
rect 10653 747 10679 749
rect 10735 747 10760 749
rect 10816 747 10841 749
rect 10897 747 10922 749
rect 10978 747 11003 749
rect 11059 747 11084 749
rect 11140 747 11149 749
tri 11149 747 11151 749 nw
tri 12099 747 12101 749 ne
rect 12101 747 12110 749
rect 12166 747 12192 749
rect 12248 747 12274 749
rect 12330 747 12356 749
rect 12412 747 12438 749
rect 12494 747 12520 749
rect 12576 747 12601 749
rect 12657 747 12682 749
rect 12738 747 12763 749
rect 12819 747 12844 749
rect 12900 747 12925 749
rect 12981 747 12990 749
tri 12990 747 12992 749 nw
tri 16742 747 16744 749 ne
rect 16744 747 16753 749
rect 16809 747 16835 749
rect 16891 747 16917 749
rect 16973 747 16999 749
rect 17055 747 17081 749
rect 17137 747 17163 749
rect 17219 747 17244 749
rect 17300 747 17325 749
rect 17381 747 17406 749
rect 17462 747 17487 749
rect 17543 747 17568 749
rect 17624 747 17633 749
tri 17633 747 17635 749 nw
tri 18583 747 18585 749 ne
rect 18585 747 18594 749
rect 18650 747 18676 749
rect 18732 747 18758 749
rect 18814 747 18840 749
rect 18896 747 18922 749
rect 18978 747 19004 749
rect 19060 747 19085 749
rect 19141 747 19166 749
rect 19222 747 19247 749
rect 19303 747 19328 749
rect 19384 747 19409 749
rect 19465 747 19474 749
tri 19474 747 19476 749 nw
rect 22236 714 22288 720
rect 22430 1803 23308 2063
rect 22430 1751 22439 1803
rect 22491 1751 22507 1803
rect 22559 1751 22575 1803
rect 22627 1751 22643 1803
rect 22695 1751 22711 1803
rect 22763 1751 22779 1803
rect 22831 1751 22847 1803
rect 22899 1751 22915 1803
rect 22967 1751 22982 1803
rect 23034 1751 23049 1803
rect 23101 1751 23116 1803
rect 23168 1751 23183 1803
rect 23235 1751 23250 1803
rect 23302 1751 23308 1803
rect 22430 1491 23308 1751
rect 22430 1439 22439 1491
rect 22491 1439 22507 1491
rect 22559 1439 22575 1491
rect 22627 1439 22643 1491
rect 22695 1439 22711 1491
rect 22763 1439 22779 1491
rect 22831 1439 22847 1491
rect 22899 1439 22915 1491
rect 22967 1439 22982 1491
rect 23034 1439 23049 1491
rect 23101 1439 23116 1491
rect 23168 1439 23183 1491
rect 23235 1439 23250 1491
rect 23302 1439 23308 1491
rect 22430 1179 23308 1439
rect 22430 1127 22439 1179
rect 22491 1127 22507 1179
rect 22559 1127 22575 1179
rect 22627 1127 22643 1179
rect 22695 1127 22711 1179
rect 22763 1127 22779 1179
rect 22831 1127 22847 1179
rect 22899 1127 22915 1179
rect 22967 1127 22982 1179
rect 23034 1127 23049 1179
rect 23101 1127 23116 1179
rect 23168 1127 23183 1179
rect 23235 1127 23250 1179
rect 23302 1127 23308 1179
rect 22430 867 23308 1127
rect 22430 815 22439 867
rect 22491 815 22507 867
rect 22559 815 22575 867
rect 22627 815 22643 867
rect 22695 815 22711 867
rect 22763 815 22779 867
rect 22831 815 22847 867
rect 22899 815 22915 867
rect 22967 815 22982 867
rect 23034 815 23049 867
rect 23101 815 23116 867
rect 23168 815 23183 867
rect 23235 815 23250 867
rect 23302 815 23308 867
tri 2348 671 2350 673 se
rect 2350 671 2359 673
rect 2415 671 2476 673
rect 2532 671 2592 673
rect 2648 671 2657 673
tri 2657 671 2659 673 sw
rect 1539 619 1545 671
rect 1597 619 1610 671
rect 1662 619 1675 671
rect 1727 619 1740 671
rect 1792 619 1805 671
rect 1857 619 1870 671
rect 1922 619 1935 671
rect 1987 619 2000 671
rect 2052 619 2065 671
rect 2117 619 2130 671
rect 2182 619 2195 671
rect 2247 619 2260 671
rect 2312 619 2325 671
rect 2442 619 2455 671
rect 2572 619 2585 671
rect 2648 619 2650 671
rect 2702 619 2715 671
rect 2767 619 2780 671
rect 2832 619 2845 671
rect 2897 619 2910 671
rect 2962 619 2975 671
rect 3027 619 3040 671
rect 3092 619 3105 671
rect 3157 619 3170 671
rect 3222 619 3235 671
rect 3287 619 3300 671
rect 3352 619 3365 671
rect 3417 619 3430 671
rect 3482 619 3495 671
rect 3547 619 3560 671
rect 3612 619 3625 671
rect 3677 619 3690 671
rect 3742 619 3755 671
rect 3807 619 3820 671
rect 3872 619 3885 671
rect 3937 619 3950 671
rect 4002 619 4015 671
rect 4067 619 4080 671
rect 4132 619 4144 671
rect 4196 619 4208 671
rect 4260 619 4272 671
rect 4324 619 4336 671
rect 4388 619 4400 671
rect 4452 619 4464 671
rect 4516 619 4528 671
rect 4580 619 4592 671
rect 4644 619 4656 671
rect 4708 619 4720 671
rect 4772 619 4784 671
rect 4836 619 4848 671
rect 4900 619 4912 671
rect 4964 619 4976 671
rect 5028 619 5040 671
rect 5092 619 5104 671
rect 5156 619 5168 671
rect 5220 619 5232 671
rect 5284 619 5296 671
rect 5348 619 5360 671
rect 5412 619 5424 671
rect 5476 619 5488 671
rect 5540 619 5552 671
rect 5604 619 5616 671
rect 5668 619 5680 671
rect 5732 619 5744 671
rect 5796 619 5808 671
rect 5860 619 5872 671
rect 5924 619 5936 671
rect 5988 619 6000 671
rect 6052 619 6064 671
rect 6116 619 6122 671
rect 22430 661 23308 815
rect 23401 1907 23407 1959
rect 23459 1907 23478 1959
rect 23530 1907 23549 1959
rect 23601 1907 23620 1959
rect 23672 1907 23691 1959
rect 23743 1907 23762 1959
rect 23814 1907 23833 1959
rect 23885 1907 23904 1959
rect 23956 1907 23975 1959
rect 24027 1907 24046 1959
rect 24098 1907 24104 1959
rect 23401 1647 24104 1907
rect 23401 1595 23407 1647
rect 23459 1595 23478 1647
rect 23530 1595 23549 1647
rect 23601 1595 23620 1647
rect 23672 1595 23691 1647
rect 23743 1595 23762 1647
rect 23814 1595 23833 1647
rect 23885 1595 23904 1647
rect 23956 1595 23975 1647
rect 24027 1595 24046 1647
rect 24098 1595 24104 1647
rect 23401 1335 24104 1595
rect 23401 1283 23407 1335
rect 23459 1283 23478 1335
rect 23530 1283 23549 1335
rect 23601 1283 23620 1335
rect 23672 1283 23691 1335
rect 23743 1283 23762 1335
rect 23814 1283 23833 1335
rect 23885 1283 23904 1335
rect 23956 1283 23975 1335
rect 24027 1283 24046 1335
rect 24098 1283 24104 1335
rect 23401 1022 24104 1283
rect 23401 970 23407 1022
rect 23459 970 23478 1022
rect 23530 970 23549 1022
rect 23601 970 23620 1022
rect 23672 970 23691 1022
rect 23743 970 23762 1022
rect 23814 970 23833 1022
rect 23885 970 23904 1022
rect 23956 970 23975 1022
rect 24027 970 24046 1022
rect 24098 970 24104 1022
rect 23401 711 24104 970
rect 23401 659 23407 711
rect 23459 659 23478 711
rect 23530 659 23549 711
rect 23601 659 23620 711
rect 23672 659 23691 711
rect 23743 659 23762 711
rect 23814 659 23833 711
rect 23885 659 23904 711
rect 23956 659 23975 711
rect 24027 659 24046 711
rect 24098 659 24104 711
rect 7714 645 7723 647
rect 7779 645 7806 647
rect 7862 645 7888 647
rect 7944 645 7970 647
rect 8026 645 8052 647
rect 8108 645 8117 647
rect 8645 645 8654 647
rect 8710 645 8737 647
rect 8793 645 8819 647
rect 8875 645 8901 647
rect 8957 645 8983 647
rect 9039 645 9048 647
rect 14198 645 14207 647
rect 14263 645 14290 647
rect 14346 645 14372 647
rect 14428 645 14454 647
rect 14510 645 14536 647
rect 14592 645 14601 647
tri 2348 617 2350 619 ne
rect 2350 617 2359 619
rect 2415 617 2476 619
rect 2532 617 2592 619
rect 2648 617 2657 619
tri 2657 617 2659 619 nw
rect 7610 593 7616 645
rect 7668 593 7681 645
rect 7798 593 7806 645
rect 7863 593 7876 645
rect 8123 593 8136 645
rect 8188 593 8201 645
rect 8253 593 8266 645
rect 8318 593 8331 645
rect 8383 593 8396 645
rect 8448 593 8461 645
rect 8513 593 8526 645
rect 8578 593 8591 645
rect 8643 593 8654 645
rect 8710 593 8721 645
rect 8968 593 8981 645
rect 9039 593 9046 645
rect 9098 593 9111 645
rect 9163 593 9176 645
rect 9228 593 9241 645
rect 9293 593 9306 645
rect 9358 593 9371 645
rect 9423 593 9436 645
rect 9488 593 9501 645
rect 9553 593 9566 645
rect 9618 593 9631 645
rect 9683 593 9696 645
rect 9748 593 9761 645
rect 9813 593 9826 645
rect 9878 593 9891 645
rect 9943 593 9956 645
rect 10008 593 10021 645
rect 10073 593 10086 645
rect 10138 593 10151 645
rect 10203 593 10216 645
rect 10268 593 10281 645
rect 10333 593 10346 645
rect 10398 593 10411 645
rect 10463 593 10476 645
rect 10528 593 10541 645
rect 10593 593 10606 645
rect 10658 593 10671 645
rect 10723 593 10736 645
rect 10788 593 10800 645
rect 10852 593 10864 645
rect 10916 593 10928 645
rect 10980 593 10992 645
rect 11044 593 11056 645
rect 11108 593 11120 645
rect 11172 593 11184 645
rect 11236 593 11248 645
rect 11300 593 11312 645
rect 11364 593 11376 645
rect 11428 593 11440 645
rect 11492 593 11504 645
rect 11556 593 11568 645
rect 11620 593 11632 645
rect 11684 593 11696 645
rect 11748 593 11760 645
rect 11812 593 11824 645
rect 11876 593 11882 645
rect 12016 593 12022 645
rect 12074 593 12087 645
rect 12139 593 12152 645
rect 12204 593 12217 645
rect 12269 593 12282 645
rect 12334 593 12347 645
rect 12399 593 12412 645
rect 12464 593 12477 645
rect 12529 593 12542 645
rect 12594 593 12607 645
rect 12659 593 12672 645
rect 12724 593 12737 645
rect 12789 593 12802 645
rect 12854 593 12867 645
rect 12919 593 12932 645
rect 12984 593 12997 645
rect 13049 593 13062 645
rect 13114 593 13127 645
rect 13179 593 13192 645
rect 13244 593 13257 645
rect 13309 593 13322 645
rect 13374 593 13387 645
rect 13439 593 13452 645
rect 13504 593 13517 645
rect 13569 593 13582 645
rect 13634 593 13647 645
rect 13699 593 13712 645
rect 13764 593 13777 645
rect 13829 593 13842 645
rect 13894 593 13907 645
rect 13959 593 13972 645
rect 14024 593 14037 645
rect 14089 593 14102 645
rect 14154 593 14167 645
rect 14284 593 14290 645
rect 14349 593 14362 645
rect 14609 593 14622 645
rect 14674 593 14687 645
rect 14739 593 14752 645
rect 14804 593 14817 645
rect 14869 593 14882 645
rect 14934 593 14947 645
rect 14999 593 15012 645
rect 15064 593 15077 645
rect 7714 591 7723 593
rect 7779 591 7806 593
rect 7862 591 7888 593
rect 7944 591 7970 593
rect 8026 591 8052 593
rect 8108 591 8117 593
rect 8645 591 8654 593
rect 8710 591 8737 593
rect 8793 591 8819 593
rect 8875 591 8901 593
rect 8957 591 8983 593
rect 9039 591 9048 593
rect 14198 591 14207 593
rect 14263 591 14290 593
rect 14346 591 14372 593
rect 14428 591 14454 593
rect 14510 591 14536 593
rect 14592 591 14601 593
rect 15129 591 15138 647
rect 15194 645 15221 647
rect 15277 645 15303 647
rect 15359 645 15385 647
rect 15441 645 15467 647
rect 15523 645 15532 647
rect 20767 645 20776 647
rect 20832 645 20858 647
rect 20914 645 20939 647
rect 20995 645 21020 647
rect 21076 645 21085 647
rect 15194 593 15206 645
rect 15450 593 15462 645
rect 15523 593 15526 645
rect 15578 593 15590 645
rect 15642 593 15654 645
rect 15706 593 15718 645
rect 15770 593 15782 645
rect 15834 593 15846 645
rect 15898 593 15910 645
rect 15962 593 15974 645
rect 16026 593 16038 645
rect 16090 593 16102 645
rect 16154 593 16166 645
rect 16218 593 16230 645
rect 16282 593 16294 645
rect 16346 593 16358 645
rect 16410 593 16422 645
rect 16474 593 16486 645
rect 16538 593 16550 645
rect 16602 593 16614 645
rect 16666 593 16678 645
rect 16730 593 16742 645
rect 16794 593 16806 645
rect 16858 593 16870 645
rect 16922 593 16934 645
rect 16986 593 16998 645
rect 17050 593 17062 645
rect 17114 593 17126 645
rect 17178 593 17190 645
rect 17242 593 17254 645
rect 17306 593 17318 645
rect 17370 593 17382 645
rect 17434 593 17446 645
rect 17498 593 17510 645
rect 17562 593 17574 645
rect 17626 593 17638 645
rect 17690 593 17702 645
rect 17754 593 17766 645
rect 17818 593 17830 645
rect 17882 593 17894 645
rect 17946 593 17958 645
rect 18010 593 18022 645
rect 18074 593 18086 645
rect 18138 593 18150 645
rect 18202 593 18214 645
rect 18266 593 18278 645
rect 18330 593 18342 645
rect 18394 593 18406 645
rect 18458 593 18470 645
rect 18522 593 18534 645
rect 18586 593 18598 645
rect 18650 593 18662 645
rect 18714 593 18726 645
rect 18778 593 18790 645
rect 18842 593 18854 645
rect 18906 593 18918 645
rect 18970 593 18982 645
rect 19034 593 19046 645
rect 19098 593 19110 645
rect 19162 593 19174 645
rect 19226 593 19238 645
rect 19290 593 19302 645
rect 19354 593 19366 645
rect 19418 593 19430 645
rect 19482 593 19494 645
rect 19546 593 19558 645
rect 19610 593 19622 645
rect 19674 593 19686 645
rect 19738 593 19750 645
rect 19802 593 19814 645
rect 19866 593 19878 645
rect 19930 593 19942 645
rect 19994 593 20006 645
rect 20058 593 20070 645
rect 20122 593 20134 645
rect 20186 593 20198 645
rect 20250 593 20262 645
rect 20314 593 20326 645
rect 20378 593 20390 645
rect 20442 593 20454 645
rect 20506 593 20518 645
rect 20570 593 20582 645
rect 20634 593 20646 645
rect 20698 593 20710 645
rect 20762 593 20774 645
rect 20832 593 20838 645
rect 21018 593 21020 645
rect 21082 593 21094 645
rect 21146 593 21158 645
rect 21210 593 21222 645
rect 21274 593 21286 645
rect 21338 593 21350 645
rect 21402 593 21414 645
rect 21466 593 21478 645
rect 21530 593 21542 645
rect 21594 593 21606 645
rect 21658 593 21670 645
rect 21722 593 21734 645
rect 21786 593 21798 645
rect 21850 593 21862 645
rect 21914 593 21926 645
rect 21978 593 21984 645
rect 15194 591 15221 593
rect 15277 591 15303 593
rect 15359 591 15385 593
rect 15441 591 15467 593
rect 15523 591 15532 593
rect 20767 591 20776 593
rect 20832 591 20858 593
rect 20914 591 20939 593
rect 20995 591 21020 593
rect 21076 591 21085 593
rect 23401 525 24104 659
rect 20688 473 20694 525
rect 20746 473 20760 525
rect 20812 503 20826 525
rect 20878 503 20892 525
rect 20944 503 20957 525
rect 21009 503 21022 525
rect 21074 503 21080 525
rect 21009 473 21019 503
rect 20688 461 20776 473
rect 20832 461 20857 473
rect 20913 461 20938 473
rect 20994 461 21019 473
rect 20688 409 20694 461
rect 20746 409 20760 461
rect 21009 447 21019 461
rect 21075 447 21084 503
rect 20812 423 20826 447
rect 20878 423 20892 447
rect 20944 423 20957 447
rect 21009 423 21022 447
rect 21074 423 21084 447
rect 21009 409 21019 423
rect 20688 397 20776 409
rect 20832 397 20857 409
rect 20913 397 20938 409
rect 20994 397 21019 409
rect 20688 345 20694 397
rect 20746 345 20760 397
rect 21009 367 21019 397
rect 21075 367 21084 423
rect 23401 473 23407 525
rect 23459 473 23478 525
rect 23530 473 23549 525
rect 23601 473 23620 525
rect 23672 473 23691 525
rect 23743 473 23761 525
rect 23813 473 23831 525
rect 23883 473 23901 525
rect 23953 473 23971 525
rect 24023 473 24041 525
rect 24093 473 24104 525
rect 23401 461 24104 473
rect 23401 409 23407 461
rect 23459 409 23478 461
rect 23530 409 23549 461
rect 23601 409 23620 461
rect 23672 409 23691 461
rect 23743 409 23761 461
rect 23813 409 23831 461
rect 23883 409 23901 461
rect 23953 409 23971 461
rect 24023 409 24041 461
rect 24093 409 24104 461
rect 23401 397 24104 409
rect 20812 345 20826 367
rect 20878 345 20892 367
rect 20944 345 20957 367
rect 21009 345 21022 367
rect 21074 345 21080 367
rect 23401 345 23407 397
rect 23459 345 23478 397
rect 23530 345 23549 397
rect 23601 345 23620 397
rect 23672 345 23691 397
rect 23743 345 23761 397
rect 23813 345 23831 397
rect 23883 345 23901 397
rect 23953 345 23971 397
rect 24023 345 24041 397
rect 24093 351 24104 397
rect 24093 345 24099 351
<< via2 >>
rect 18590 2972 18646 3028
rect 18672 2972 18728 3028
rect 18754 2972 18810 3028
rect 18836 2972 18892 3028
rect 18918 2972 18974 3028
rect 19000 2972 19056 3028
rect 19082 2972 19138 3028
rect 19164 2972 19220 3028
rect 19247 2972 19303 3028
rect 19330 2972 19386 3028
rect 19413 2972 19469 3028
rect 18590 2838 18646 2894
rect 18672 2838 18728 2894
rect 18754 2838 18810 2894
rect 18836 2838 18892 2894
rect 18918 2838 18974 2894
rect 19000 2838 19056 2894
rect 19082 2838 19138 2894
rect 19164 2838 19220 2894
rect 19247 2838 19303 2894
rect 19330 2838 19386 2894
rect 19413 2838 19469 2894
rect 7723 1269 7779 1271
rect 7806 1269 7862 1271
rect 7888 1269 7944 1271
rect 7970 1269 8026 1271
rect 8052 1269 8108 1271
rect 8654 1269 8710 1271
rect 8737 1269 8793 1271
rect 8819 1269 8875 1271
rect 8901 1269 8957 1271
rect 8983 1269 9039 1271
rect 14211 1270 14267 1271
rect 14294 1270 14350 1271
rect 14376 1270 14432 1271
rect 14458 1270 14514 1271
rect 14540 1270 14596 1271
rect 15138 1270 15194 1271
rect 15221 1270 15277 1271
rect 15303 1270 15359 1271
rect 15385 1270 15441 1271
rect 15467 1270 15523 1271
rect 20776 1270 20832 1271
rect 20859 1270 20915 1271
rect 20942 1270 20998 1271
rect 21024 1270 21080 1271
rect 7723 1217 7733 1269
rect 7733 1217 7746 1269
rect 7746 1217 7779 1269
rect 7806 1217 7811 1269
rect 7811 1217 7862 1269
rect 7888 1217 7928 1269
rect 7928 1217 7941 1269
rect 7941 1217 7944 1269
rect 7970 1217 7993 1269
rect 7993 1217 8006 1269
rect 8006 1217 8026 1269
rect 8052 1217 8058 1269
rect 8058 1217 8071 1269
rect 8071 1217 8108 1269
rect 8654 1217 8656 1269
rect 8656 1217 8708 1269
rect 8708 1217 8710 1269
rect 8737 1217 8773 1269
rect 8773 1217 8786 1269
rect 8786 1217 8793 1269
rect 8819 1217 8838 1269
rect 8838 1217 8851 1269
rect 8851 1217 8875 1269
rect 8901 1217 8903 1269
rect 8903 1217 8916 1269
rect 8916 1217 8957 1269
rect 8983 1217 9033 1269
rect 9033 1217 9039 1269
rect 14211 1218 14261 1270
rect 14261 1218 14267 1270
rect 14294 1218 14325 1270
rect 14325 1218 14337 1270
rect 14337 1218 14350 1270
rect 14376 1218 14389 1270
rect 14389 1218 14401 1270
rect 14401 1218 14432 1270
rect 14458 1218 14465 1270
rect 14465 1218 14514 1270
rect 14540 1218 14581 1270
rect 14581 1218 14593 1270
rect 14593 1218 14596 1270
rect 15138 1218 15157 1270
rect 15157 1218 15169 1270
rect 15169 1218 15194 1270
rect 15221 1218 15233 1270
rect 15233 1218 15277 1270
rect 15303 1218 15349 1270
rect 15349 1218 15359 1270
rect 15385 1218 15413 1270
rect 15413 1218 15425 1270
rect 15425 1218 15441 1270
rect 15467 1218 15477 1270
rect 15477 1218 15489 1270
rect 15489 1218 15523 1270
rect 20776 1218 20789 1270
rect 20789 1218 20801 1270
rect 20801 1218 20832 1270
rect 20859 1218 20865 1270
rect 20865 1218 20915 1270
rect 20942 1218 20981 1270
rect 20981 1218 20993 1270
rect 20993 1218 20998 1270
rect 21024 1218 21045 1270
rect 21045 1218 21057 1270
rect 21057 1218 21080 1270
rect 7723 1215 7779 1217
rect 7806 1215 7862 1217
rect 7888 1215 7944 1217
rect 7970 1215 8026 1217
rect 8052 1215 8108 1217
rect 8654 1215 8710 1217
rect 8737 1215 8793 1217
rect 8819 1215 8875 1217
rect 8901 1215 8957 1217
rect 8983 1215 9039 1217
rect 14211 1215 14267 1218
rect 14294 1215 14350 1218
rect 14376 1215 14432 1218
rect 14458 1215 14514 1218
rect 14540 1215 14596 1218
rect 15138 1215 15194 1218
rect 15221 1215 15277 1218
rect 15303 1215 15359 1218
rect 15385 1215 15441 1218
rect 15467 1215 15523 1218
rect 20776 1215 20832 1218
rect 20859 1215 20915 1218
rect 20942 1215 20998 1218
rect 21024 1215 21080 1218
rect 10269 1113 10325 1115
rect 10351 1113 10407 1115
rect 10433 1113 10489 1115
rect 10515 1113 10571 1115
rect 10597 1113 10653 1115
rect 10679 1113 10735 1115
rect 10760 1113 10816 1115
rect 10841 1113 10897 1115
rect 10922 1113 10978 1115
rect 11003 1113 11059 1115
rect 11084 1113 11140 1115
rect 12110 1113 12166 1115
rect 12192 1113 12248 1115
rect 12274 1113 12330 1115
rect 12356 1113 12412 1115
rect 12438 1113 12494 1115
rect 12520 1113 12576 1115
rect 12601 1113 12657 1115
rect 12682 1113 12738 1115
rect 12763 1113 12819 1115
rect 12844 1113 12900 1115
rect 12925 1113 12981 1115
rect 16753 1113 16809 1115
rect 16835 1113 16891 1115
rect 16917 1113 16973 1115
rect 16999 1113 17055 1115
rect 17081 1113 17137 1115
rect 17163 1113 17219 1115
rect 17244 1113 17300 1115
rect 17325 1113 17381 1115
rect 17406 1113 17462 1115
rect 17487 1113 17543 1115
rect 17568 1113 17624 1115
rect 18594 1113 18650 1115
rect 18676 1113 18732 1115
rect 18758 1113 18814 1115
rect 18840 1113 18896 1115
rect 18922 1113 18978 1115
rect 19004 1113 19060 1115
rect 19085 1113 19141 1115
rect 19166 1113 19222 1115
rect 19247 1113 19303 1115
rect 19328 1113 19384 1115
rect 19409 1113 19465 1115
rect 10269 1061 10281 1113
rect 10281 1061 10325 1113
rect 10351 1061 10398 1113
rect 10398 1061 10407 1113
rect 10433 1061 10463 1113
rect 10463 1061 10476 1113
rect 10476 1061 10489 1113
rect 10515 1061 10528 1113
rect 10528 1061 10541 1113
rect 10541 1061 10571 1113
rect 10597 1061 10606 1113
rect 10606 1061 10653 1113
rect 10679 1061 10723 1113
rect 10723 1061 10735 1113
rect 10760 1061 10788 1113
rect 10788 1061 10800 1113
rect 10800 1061 10816 1113
rect 10841 1061 10852 1113
rect 10852 1061 10864 1113
rect 10864 1061 10897 1113
rect 10922 1061 10928 1113
rect 10928 1061 10978 1113
rect 11003 1061 11044 1113
rect 11044 1061 11056 1113
rect 11056 1061 11059 1113
rect 11084 1061 11108 1113
rect 11108 1061 11120 1113
rect 11120 1061 11140 1113
rect 12110 1061 12139 1113
rect 12139 1061 12152 1113
rect 12152 1061 12166 1113
rect 12192 1061 12204 1113
rect 12204 1061 12217 1113
rect 12217 1061 12248 1113
rect 12274 1061 12282 1113
rect 12282 1061 12330 1113
rect 12356 1061 12399 1113
rect 12399 1061 12412 1113
rect 12438 1061 12464 1113
rect 12464 1061 12477 1113
rect 12477 1061 12494 1113
rect 12520 1061 12529 1113
rect 12529 1061 12542 1113
rect 12542 1061 12576 1113
rect 12601 1061 12607 1113
rect 12607 1061 12657 1113
rect 12682 1061 12724 1113
rect 12724 1061 12737 1113
rect 12737 1061 12738 1113
rect 12763 1061 12789 1113
rect 12789 1061 12801 1113
rect 12801 1061 12819 1113
rect 12844 1061 12853 1113
rect 12853 1061 12865 1113
rect 12865 1061 12900 1113
rect 12925 1061 12929 1113
rect 12929 1061 12981 1113
rect 16753 1061 16757 1113
rect 16757 1061 16769 1113
rect 16769 1061 16809 1113
rect 16835 1061 16885 1113
rect 16885 1061 16891 1113
rect 16917 1061 16949 1113
rect 16949 1061 16961 1113
rect 16961 1061 16973 1113
rect 16999 1061 17013 1113
rect 17013 1061 17025 1113
rect 17025 1061 17055 1113
rect 17081 1061 17089 1113
rect 17089 1061 17137 1113
rect 17163 1061 17205 1113
rect 17205 1061 17217 1113
rect 17217 1061 17219 1113
rect 17244 1061 17269 1113
rect 17269 1061 17281 1113
rect 17281 1061 17300 1113
rect 17325 1061 17333 1113
rect 17333 1061 17345 1113
rect 17345 1061 17381 1113
rect 17406 1061 17409 1113
rect 17409 1061 17461 1113
rect 17461 1061 17462 1113
rect 17487 1061 17525 1113
rect 17525 1061 17537 1113
rect 17537 1061 17543 1113
rect 17568 1061 17589 1113
rect 17589 1061 17601 1113
rect 17601 1061 17624 1113
rect 18594 1061 18613 1113
rect 18613 1061 18625 1113
rect 18625 1061 18650 1113
rect 18676 1061 18677 1113
rect 18677 1061 18689 1113
rect 18689 1061 18732 1113
rect 18758 1061 18805 1113
rect 18805 1061 18814 1113
rect 18840 1061 18869 1113
rect 18869 1061 18881 1113
rect 18881 1061 18896 1113
rect 18922 1061 18933 1113
rect 18933 1061 18945 1113
rect 18945 1061 18978 1113
rect 19004 1061 19009 1113
rect 19009 1061 19060 1113
rect 19085 1061 19125 1113
rect 19125 1061 19137 1113
rect 19137 1061 19141 1113
rect 19166 1061 19189 1113
rect 19189 1061 19201 1113
rect 19201 1061 19222 1113
rect 19247 1061 19253 1113
rect 19253 1061 19265 1113
rect 19265 1061 19303 1113
rect 19328 1061 19329 1113
rect 19329 1061 19381 1113
rect 19381 1061 19384 1113
rect 19409 1061 19445 1113
rect 19445 1061 19457 1113
rect 19457 1061 19465 1113
rect 10269 1059 10325 1061
rect 10351 1059 10407 1061
rect 10433 1059 10489 1061
rect 10515 1059 10571 1061
rect 10597 1059 10653 1061
rect 10679 1059 10735 1061
rect 10760 1059 10816 1061
rect 10841 1059 10897 1061
rect 10922 1059 10978 1061
rect 11003 1059 11059 1061
rect 11084 1059 11140 1061
rect 12110 1059 12166 1061
rect 12192 1059 12248 1061
rect 12274 1059 12330 1061
rect 12356 1059 12412 1061
rect 12438 1059 12494 1061
rect 12520 1059 12576 1061
rect 12601 1059 12657 1061
rect 12682 1059 12738 1061
rect 12763 1059 12819 1061
rect 12844 1059 12900 1061
rect 12925 1059 12981 1061
rect 16753 1059 16809 1061
rect 16835 1059 16891 1061
rect 16917 1059 16973 1061
rect 16999 1059 17055 1061
rect 17081 1059 17137 1061
rect 17163 1059 17219 1061
rect 17244 1059 17300 1061
rect 17325 1059 17381 1061
rect 17406 1059 17462 1061
rect 17487 1059 17543 1061
rect 17568 1059 17624 1061
rect 18594 1059 18650 1061
rect 18676 1059 18732 1061
rect 18758 1059 18814 1061
rect 18840 1059 18896 1061
rect 18922 1059 18978 1061
rect 19004 1059 19060 1061
rect 19085 1059 19141 1061
rect 19166 1059 19222 1061
rect 19247 1059 19303 1061
rect 19328 1059 19384 1061
rect 19409 1059 19465 1061
rect 7723 957 7779 959
rect 7806 957 7862 959
rect 7888 957 7944 959
rect 7970 957 8026 959
rect 8052 957 8108 959
rect 8654 957 8710 959
rect 8737 957 8793 959
rect 8819 957 8875 959
rect 8901 957 8957 959
rect 8983 957 9039 959
rect 14207 957 14263 959
rect 14290 957 14346 959
rect 14372 957 14428 959
rect 14454 957 14510 959
rect 14536 957 14592 959
rect 15138 957 15194 959
rect 15221 957 15277 959
rect 15303 957 15359 959
rect 15385 957 15441 959
rect 15467 957 15523 959
rect 20776 957 20832 959
rect 20858 957 20914 959
rect 20939 957 20995 959
rect 21020 957 21076 959
rect 7723 905 7733 957
rect 7733 905 7746 957
rect 7746 905 7779 957
rect 7806 905 7811 957
rect 7811 905 7862 957
rect 7888 905 7928 957
rect 7928 905 7941 957
rect 7941 905 7944 957
rect 7970 905 7993 957
rect 7993 905 8006 957
rect 8006 905 8026 957
rect 8052 905 8058 957
rect 8058 905 8071 957
rect 8071 905 8108 957
rect 8654 905 8656 957
rect 8656 905 8708 957
rect 8708 905 8710 957
rect 8737 905 8773 957
rect 8773 905 8786 957
rect 8786 905 8793 957
rect 8819 905 8838 957
rect 8838 905 8851 957
rect 8851 905 8875 957
rect 8901 905 8903 957
rect 8903 905 8916 957
rect 8916 905 8957 957
rect 8983 905 9033 957
rect 9033 905 9039 957
rect 14207 905 14219 957
rect 14219 905 14232 957
rect 14232 905 14263 957
rect 14290 905 14297 957
rect 14297 905 14346 957
rect 14372 905 14414 957
rect 14414 905 14427 957
rect 14427 905 14428 957
rect 14454 905 14479 957
rect 14479 905 14492 957
rect 14492 905 14510 957
rect 14536 905 14544 957
rect 14544 905 14557 957
rect 14557 905 14592 957
rect 15138 905 15186 957
rect 15186 905 15194 957
rect 15221 905 15250 957
rect 15250 905 15262 957
rect 15262 905 15277 957
rect 15303 905 15314 957
rect 15314 905 15326 957
rect 15326 905 15359 957
rect 15385 905 15390 957
rect 15390 905 15441 957
rect 15467 905 15506 957
rect 15506 905 15518 957
rect 15518 905 15523 957
rect 20776 905 20818 957
rect 20818 905 20830 957
rect 20830 905 20832 957
rect 20858 905 20882 957
rect 20882 905 20894 957
rect 20894 905 20914 957
rect 20939 905 20946 957
rect 20946 905 20958 957
rect 20958 905 20995 957
rect 21020 905 21022 957
rect 21022 905 21074 957
rect 21074 905 21076 957
rect 7723 903 7779 905
rect 7806 903 7862 905
rect 7888 903 7944 905
rect 7970 903 8026 905
rect 8052 903 8108 905
rect 8654 903 8710 905
rect 8737 903 8793 905
rect 8819 903 8875 905
rect 8901 903 8957 905
rect 8983 903 9039 905
rect 14207 903 14263 905
rect 14290 903 14346 905
rect 14372 903 14428 905
rect 14454 903 14510 905
rect 14536 903 14592 905
rect 15138 903 15194 905
rect 15221 903 15277 905
rect 15303 903 15359 905
rect 15385 903 15441 905
rect 15467 903 15523 905
rect 20776 903 20832 905
rect 20858 903 20914 905
rect 20939 903 20995 905
rect 21020 903 21076 905
rect 5626 827 5682 829
rect 5714 827 5770 829
rect 5802 827 5858 829
rect 5890 827 5946 829
rect 5978 827 6034 829
rect 6066 827 6122 829
rect 5626 775 5668 827
rect 5668 775 5680 827
rect 5680 775 5682 827
rect 5714 775 5732 827
rect 5732 775 5744 827
rect 5744 775 5770 827
rect 5802 775 5808 827
rect 5808 775 5858 827
rect 5890 775 5924 827
rect 5924 775 5936 827
rect 5936 775 5946 827
rect 5978 775 5988 827
rect 5988 775 6000 827
rect 6000 775 6034 827
rect 6066 775 6116 827
rect 6116 775 6122 827
rect 5626 773 5682 775
rect 5714 773 5770 775
rect 5802 773 5858 775
rect 5890 773 5946 775
rect 5978 773 6034 775
rect 6066 773 6122 775
rect 6153 773 6209 829
rect 10269 801 10325 803
rect 10351 801 10407 803
rect 10433 801 10489 803
rect 10515 801 10571 803
rect 10597 801 10653 803
rect 10679 801 10735 803
rect 10760 801 10816 803
rect 10841 801 10897 803
rect 10922 801 10978 803
rect 11003 801 11059 803
rect 11084 801 11140 803
rect 12110 801 12166 803
rect 12192 801 12248 803
rect 12274 801 12330 803
rect 12356 801 12412 803
rect 12438 801 12494 803
rect 12520 801 12576 803
rect 12601 801 12657 803
rect 12682 801 12738 803
rect 12763 801 12819 803
rect 12844 801 12900 803
rect 12925 801 12981 803
rect 16753 801 16809 803
rect 16835 801 16891 803
rect 16917 801 16973 803
rect 16999 801 17055 803
rect 17081 801 17137 803
rect 17163 801 17219 803
rect 17244 801 17300 803
rect 17325 801 17381 803
rect 17406 801 17462 803
rect 17487 801 17543 803
rect 17568 801 17624 803
rect 18594 801 18650 803
rect 18676 801 18732 803
rect 18758 801 18814 803
rect 18840 801 18896 803
rect 18922 801 18978 803
rect 19004 801 19060 803
rect 19085 801 19141 803
rect 19166 801 19222 803
rect 19247 801 19303 803
rect 19328 801 19384 803
rect 19409 801 19465 803
rect 10269 749 10281 801
rect 10281 749 10325 801
rect 10351 749 10398 801
rect 10398 749 10407 801
rect 10433 749 10463 801
rect 10463 749 10476 801
rect 10476 749 10489 801
rect 10515 749 10528 801
rect 10528 749 10541 801
rect 10541 749 10571 801
rect 10597 749 10606 801
rect 10606 749 10653 801
rect 10679 749 10723 801
rect 10723 749 10735 801
rect 10760 749 10788 801
rect 10788 749 10800 801
rect 10800 749 10816 801
rect 10841 749 10852 801
rect 10852 749 10864 801
rect 10864 749 10897 801
rect 10922 749 10928 801
rect 10928 749 10978 801
rect 11003 749 11044 801
rect 11044 749 11056 801
rect 11056 749 11059 801
rect 11084 749 11108 801
rect 11108 749 11120 801
rect 11120 749 11140 801
rect 12110 749 12139 801
rect 12139 749 12152 801
rect 12152 749 12166 801
rect 12192 749 12204 801
rect 12204 749 12217 801
rect 12217 749 12248 801
rect 12274 749 12282 801
rect 12282 749 12330 801
rect 12356 749 12399 801
rect 12399 749 12412 801
rect 12438 749 12464 801
rect 12464 749 12477 801
rect 12477 749 12494 801
rect 12520 749 12529 801
rect 12529 749 12542 801
rect 12542 749 12576 801
rect 12601 749 12607 801
rect 12607 749 12657 801
rect 12682 749 12724 801
rect 12724 749 12737 801
rect 12737 749 12738 801
rect 12763 749 12789 801
rect 12789 749 12802 801
rect 12802 749 12819 801
rect 12844 749 12854 801
rect 12854 749 12867 801
rect 12867 749 12900 801
rect 12925 749 12932 801
rect 12932 749 12981 801
rect 16753 749 16777 801
rect 16777 749 16789 801
rect 16789 749 16809 801
rect 16835 749 16841 801
rect 16841 749 16853 801
rect 16853 749 16891 801
rect 16917 749 16969 801
rect 16969 749 16973 801
rect 16999 749 17033 801
rect 17033 749 17045 801
rect 17045 749 17055 801
rect 17081 749 17097 801
rect 17097 749 17109 801
rect 17109 749 17137 801
rect 17163 749 17173 801
rect 17173 749 17219 801
rect 17244 749 17289 801
rect 17289 749 17300 801
rect 17325 749 17353 801
rect 17353 749 17365 801
rect 17365 749 17381 801
rect 17406 749 17417 801
rect 17417 749 17429 801
rect 17429 749 17462 801
rect 17487 749 17493 801
rect 17493 749 17543 801
rect 17568 749 17609 801
rect 17609 749 17621 801
rect 17621 749 17624 801
rect 18594 749 18633 801
rect 18633 749 18645 801
rect 18645 749 18650 801
rect 18676 749 18697 801
rect 18697 749 18709 801
rect 18709 749 18732 801
rect 18758 749 18761 801
rect 18761 749 18773 801
rect 18773 749 18814 801
rect 18840 749 18889 801
rect 18889 749 18896 801
rect 18922 749 18953 801
rect 18953 749 18965 801
rect 18965 749 18978 801
rect 19004 749 19017 801
rect 19017 749 19029 801
rect 19029 749 19060 801
rect 19085 749 19093 801
rect 19093 749 19141 801
rect 19166 749 19209 801
rect 19209 749 19221 801
rect 19221 749 19222 801
rect 19247 749 19273 801
rect 19273 749 19285 801
rect 19285 749 19303 801
rect 19328 749 19337 801
rect 19337 749 19349 801
rect 19349 749 19384 801
rect 19409 749 19413 801
rect 19413 749 19465 801
rect 10269 747 10325 749
rect 10351 747 10407 749
rect 10433 747 10489 749
rect 10515 747 10571 749
rect 10597 747 10653 749
rect 10679 747 10735 749
rect 10760 747 10816 749
rect 10841 747 10897 749
rect 10922 747 10978 749
rect 11003 747 11059 749
rect 11084 747 11140 749
rect 12110 747 12166 749
rect 12192 747 12248 749
rect 12274 747 12330 749
rect 12356 747 12412 749
rect 12438 747 12494 749
rect 12520 747 12576 749
rect 12601 747 12657 749
rect 12682 747 12738 749
rect 12763 747 12819 749
rect 12844 747 12900 749
rect 12925 747 12981 749
rect 16753 747 16809 749
rect 16835 747 16891 749
rect 16917 747 16973 749
rect 16999 747 17055 749
rect 17081 747 17137 749
rect 17163 747 17219 749
rect 17244 747 17300 749
rect 17325 747 17381 749
rect 17406 747 17462 749
rect 17487 747 17543 749
rect 17568 747 17624 749
rect 18594 747 18650 749
rect 18676 747 18732 749
rect 18758 747 18814 749
rect 18840 747 18896 749
rect 18922 747 18978 749
rect 19004 747 19060 749
rect 19085 747 19141 749
rect 19166 747 19222 749
rect 19247 747 19303 749
rect 19328 747 19384 749
rect 19409 747 19465 749
rect 2359 671 2415 673
rect 2476 671 2532 673
rect 2592 671 2648 673
rect 2359 619 2377 671
rect 2377 619 2390 671
rect 2390 619 2415 671
rect 2476 619 2507 671
rect 2507 619 2520 671
rect 2520 619 2532 671
rect 2592 619 2637 671
rect 2637 619 2648 671
rect 7723 645 7779 647
rect 7806 645 7862 647
rect 7888 645 7944 647
rect 7970 645 8026 647
rect 8052 645 8108 647
rect 8654 645 8710 647
rect 8737 645 8793 647
rect 8819 645 8875 647
rect 8901 645 8957 647
rect 8983 645 9039 647
rect 14207 645 14263 647
rect 14290 645 14346 647
rect 14372 645 14428 647
rect 14454 645 14510 647
rect 14536 645 14592 647
rect 2359 617 2415 619
rect 2476 617 2532 619
rect 2592 617 2648 619
rect 7723 593 7733 645
rect 7733 593 7746 645
rect 7746 593 7779 645
rect 7806 593 7811 645
rect 7811 593 7862 645
rect 7888 593 7928 645
rect 7928 593 7941 645
rect 7941 593 7944 645
rect 7970 593 7993 645
rect 7993 593 8006 645
rect 8006 593 8026 645
rect 8052 593 8058 645
rect 8058 593 8071 645
rect 8071 593 8108 645
rect 8654 593 8656 645
rect 8656 593 8708 645
rect 8708 593 8710 645
rect 8737 593 8773 645
rect 8773 593 8786 645
rect 8786 593 8793 645
rect 8819 593 8838 645
rect 8838 593 8851 645
rect 8851 593 8875 645
rect 8901 593 8903 645
rect 8903 593 8916 645
rect 8916 593 8957 645
rect 8983 593 9033 645
rect 9033 593 9039 645
rect 14207 593 14219 645
rect 14219 593 14232 645
rect 14232 593 14263 645
rect 14290 593 14297 645
rect 14297 593 14346 645
rect 14372 593 14414 645
rect 14414 593 14427 645
rect 14427 593 14428 645
rect 14454 593 14479 645
rect 14479 593 14492 645
rect 14492 593 14510 645
rect 14536 593 14544 645
rect 14544 593 14557 645
rect 14557 593 14592 645
rect 7723 591 7779 593
rect 7806 591 7862 593
rect 7888 591 7944 593
rect 7970 591 8026 593
rect 8052 591 8108 593
rect 8654 591 8710 593
rect 8737 591 8793 593
rect 8819 591 8875 593
rect 8901 591 8957 593
rect 8983 591 9039 593
rect 14207 591 14263 593
rect 14290 591 14346 593
rect 14372 591 14428 593
rect 14454 591 14510 593
rect 14536 591 14592 593
rect 15138 645 15194 647
rect 15221 645 15277 647
rect 15303 645 15359 647
rect 15385 645 15441 647
rect 15467 645 15523 647
rect 20776 645 20832 647
rect 20858 645 20914 647
rect 20939 645 20995 647
rect 21020 645 21076 647
rect 15138 593 15142 645
rect 15142 593 15194 645
rect 15221 593 15258 645
rect 15258 593 15270 645
rect 15270 593 15277 645
rect 15303 593 15322 645
rect 15322 593 15334 645
rect 15334 593 15359 645
rect 15385 593 15386 645
rect 15386 593 15398 645
rect 15398 593 15441 645
rect 15467 593 15514 645
rect 15514 593 15523 645
rect 20776 593 20826 645
rect 20826 593 20832 645
rect 20858 593 20890 645
rect 20890 593 20902 645
rect 20902 593 20914 645
rect 20939 593 20954 645
rect 20954 593 20966 645
rect 20966 593 20995 645
rect 21020 593 21030 645
rect 21030 593 21076 645
rect 15138 591 15194 593
rect 15221 591 15277 593
rect 15303 591 15359 593
rect 15385 591 15441 593
rect 15467 591 15523 593
rect 20776 591 20832 593
rect 20858 591 20914 593
rect 20939 591 20995 593
rect 21020 591 21076 593
rect 20776 473 20812 503
rect 20812 473 20826 503
rect 20826 473 20832 503
rect 20857 473 20878 503
rect 20878 473 20892 503
rect 20892 473 20913 503
rect 20938 473 20944 503
rect 20944 473 20957 503
rect 20957 473 20994 503
rect 21019 473 21022 503
rect 21022 473 21074 503
rect 21074 473 21075 503
rect 20776 461 20832 473
rect 20857 461 20913 473
rect 20938 461 20994 473
rect 21019 461 21075 473
rect 20776 447 20812 461
rect 20812 447 20826 461
rect 20826 447 20832 461
rect 20857 447 20878 461
rect 20878 447 20892 461
rect 20892 447 20913 461
rect 20938 447 20944 461
rect 20944 447 20957 461
rect 20957 447 20994 461
rect 21019 447 21022 461
rect 21022 447 21074 461
rect 21074 447 21075 461
rect 20776 409 20812 423
rect 20812 409 20826 423
rect 20826 409 20832 423
rect 20857 409 20878 423
rect 20878 409 20892 423
rect 20892 409 20913 423
rect 20938 409 20944 423
rect 20944 409 20957 423
rect 20957 409 20994 423
rect 21019 409 21022 423
rect 21022 409 21074 423
rect 21074 409 21075 423
rect 20776 397 20832 409
rect 20857 397 20913 409
rect 20938 397 20994 409
rect 21019 397 21075 409
rect 20776 367 20812 397
rect 20812 367 20826 397
rect 20826 367 20832 397
rect 20857 367 20878 397
rect 20878 367 20892 397
rect 20892 367 20913 397
rect 20938 367 20944 397
rect 20944 367 20957 397
rect 20957 367 20994 397
rect 21019 367 21022 397
rect 21022 367 21074 397
rect 21074 367 21075 397
<< metal3 >>
rect 18585 3028 19474 3857
rect 18585 2972 18590 3028
rect 18646 2972 18672 3028
rect 18728 2972 18754 3028
rect 18810 2972 18836 3028
rect 18892 2972 18918 3028
rect 18974 2972 19000 3028
rect 19056 2972 19082 3028
rect 19138 2972 19164 3028
rect 19220 2972 19247 3028
rect 19303 2972 19330 3028
rect 19386 2972 19413 3028
rect 19469 2972 19474 3028
rect 18585 2894 19474 2972
rect 18585 2838 18590 2894
rect 18646 2838 18672 2894
rect 18728 2838 18754 2894
rect 18810 2838 18836 2894
rect 18892 2838 18918 2894
rect 18974 2838 19000 2894
rect 19056 2838 19082 2894
rect 19138 2838 19164 2894
rect 19220 2838 19247 2894
rect 19303 2838 19330 2894
rect 19386 2838 19413 2894
rect 19469 2838 19474 2894
rect 7718 1271 8113 1276
rect 7718 1215 7723 1271
rect 7779 1215 7806 1271
rect 7862 1215 7888 1271
rect 7944 1215 7970 1271
rect 8026 1215 8052 1271
rect 8108 1215 8113 1271
rect 7718 1210 8113 1215
rect 8649 1271 9044 1276
rect 8649 1215 8654 1271
rect 8710 1215 8737 1271
rect 8793 1215 8819 1271
rect 8875 1215 8901 1271
rect 8957 1215 8983 1271
rect 9039 1215 9044 1271
rect 8649 1210 9044 1215
rect 14206 1271 14601 1276
rect 14206 1215 14211 1271
rect 14267 1215 14294 1271
rect 14350 1215 14376 1271
rect 14432 1215 14458 1271
rect 14514 1215 14540 1271
rect 14596 1215 14601 1271
rect 14206 1210 14601 1215
rect 15133 1271 15528 1276
rect 15133 1215 15138 1271
rect 15194 1215 15221 1271
rect 15277 1215 15303 1271
rect 15359 1215 15385 1271
rect 15441 1215 15467 1271
rect 15523 1215 15528 1271
rect 15133 1210 15528 1215
rect 10264 1115 11145 1120
rect 10264 1059 10269 1115
rect 10325 1059 10351 1115
rect 10407 1059 10433 1115
rect 10489 1059 10515 1115
rect 10571 1059 10597 1115
rect 10653 1059 10679 1115
rect 10735 1059 10760 1115
rect 10816 1059 10841 1115
rect 10897 1059 10922 1115
rect 10978 1059 11003 1115
rect 11059 1059 11084 1115
rect 11140 1059 11145 1115
rect 10264 1054 11145 1059
rect 12105 1115 12986 1120
rect 12105 1059 12110 1115
rect 12166 1059 12192 1115
rect 12248 1059 12274 1115
rect 12330 1059 12356 1115
rect 12412 1059 12438 1115
rect 12494 1059 12520 1115
rect 12576 1059 12601 1115
rect 12657 1059 12682 1115
rect 12738 1059 12763 1115
rect 12819 1059 12844 1115
rect 12900 1059 12925 1115
rect 12981 1059 12986 1115
rect 12105 1054 12986 1059
rect 16748 1115 17629 1120
rect 16748 1059 16753 1115
rect 16809 1059 16835 1115
rect 16891 1059 16917 1115
rect 16973 1059 16999 1115
rect 17055 1059 17081 1115
rect 17137 1059 17163 1115
rect 17219 1059 17244 1115
rect 17300 1059 17325 1115
rect 17381 1059 17406 1115
rect 17462 1059 17487 1115
rect 17543 1059 17568 1115
rect 17624 1059 17629 1115
rect 16748 1054 17629 1059
rect 18585 1115 19474 2838
rect 18585 1059 18594 1115
rect 18650 1059 18676 1115
rect 18732 1059 18758 1115
rect 18814 1059 18840 1115
rect 18896 1059 18922 1115
rect 18978 1059 19004 1115
rect 19060 1059 19085 1115
rect 19141 1059 19166 1115
rect 19222 1059 19247 1115
rect 19303 1059 19328 1115
rect 19384 1059 19409 1115
rect 19465 1059 19474 1115
rect 7718 959 8113 964
rect 7718 903 7723 959
rect 7779 903 7806 959
rect 7862 903 7888 959
rect 7944 903 7970 959
rect 8026 903 8052 959
rect 8108 903 8113 959
rect 7718 898 8113 903
rect 8649 959 9044 964
rect 8649 903 8654 959
rect 8710 903 8737 959
rect 8793 903 8819 959
rect 8875 903 8901 959
rect 8957 903 8983 959
rect 9039 903 9044 959
rect 8649 898 9044 903
rect 14202 959 14597 964
rect 14202 903 14207 959
rect 14263 903 14290 959
rect 14346 903 14372 959
rect 14428 903 14454 959
rect 14510 903 14536 959
rect 14592 903 14597 959
rect 14202 898 14597 903
rect 15133 959 15528 964
rect 15133 903 15138 959
rect 15194 903 15221 959
rect 15277 903 15303 959
rect 15359 903 15385 959
rect 15441 903 15467 959
rect 15523 903 15528 959
rect 15133 898 15528 903
rect 5621 829 6214 834
rect 5621 773 5626 829
rect 5682 773 5714 829
rect 5770 773 5802 829
rect 5858 773 5890 829
rect 5946 773 5978 829
rect 6034 773 6066 829
rect 6122 773 6153 829
rect 6209 773 6214 829
rect 5621 768 6214 773
rect 10264 803 11145 808
rect 10264 747 10269 803
rect 10325 747 10351 803
rect 10407 747 10433 803
rect 10489 747 10515 803
rect 10571 747 10597 803
rect 10653 747 10679 803
rect 10735 747 10760 803
rect 10816 747 10841 803
rect 10897 747 10922 803
rect 10978 747 11003 803
rect 11059 747 11084 803
rect 11140 747 11145 803
rect 10264 742 11145 747
rect 12105 803 12986 808
rect 12105 747 12110 803
rect 12166 747 12192 803
rect 12248 747 12274 803
rect 12330 747 12356 803
rect 12412 747 12438 803
rect 12494 747 12520 803
rect 12576 747 12601 803
rect 12657 747 12682 803
rect 12738 747 12763 803
rect 12819 747 12844 803
rect 12900 747 12925 803
rect 12981 747 12986 803
rect 12105 742 12986 747
rect 16748 803 17629 808
rect 16748 747 16753 803
rect 16809 747 16835 803
rect 16891 747 16917 803
rect 16973 747 16999 803
rect 17055 747 17081 803
rect 17137 747 17163 803
rect 17219 747 17244 803
rect 17300 747 17325 803
rect 17381 747 17406 803
rect 17462 747 17487 803
rect 17543 747 17568 803
rect 17624 747 17629 803
rect 16748 742 17629 747
rect 18585 803 19474 1059
rect 18585 747 18594 803
rect 18650 747 18676 803
rect 18732 747 18758 803
rect 18814 747 18840 803
rect 18896 747 18922 803
rect 18978 747 19004 803
rect 19060 747 19085 803
rect 19141 747 19166 803
rect 19222 747 19247 803
rect 19303 747 19328 803
rect 19384 747 19409 803
rect 19465 747 19474 803
rect 2354 673 2653 678
rect 2354 617 2359 673
rect 2415 617 2476 673
rect 2532 617 2592 673
rect 2648 617 2653 673
rect 2354 612 2653 617
rect 7718 647 8113 652
rect 7718 591 7723 647
rect 7779 591 7806 647
rect 7862 591 7888 647
rect 7944 591 7970 647
rect 8026 591 8052 647
rect 8108 591 8113 647
rect 7718 586 8113 591
rect 8649 647 9044 652
rect 8649 591 8654 647
rect 8710 591 8737 647
rect 8793 591 8819 647
rect 8875 591 8901 647
rect 8957 591 8983 647
rect 9039 591 9044 647
rect 8649 586 9044 591
rect 14202 647 14597 652
rect 14202 591 14207 647
rect 14263 591 14290 647
rect 14346 591 14372 647
rect 14428 591 14454 647
rect 14510 591 14536 647
rect 14592 591 14597 647
rect 14202 586 14597 591
rect 15133 647 15528 652
rect 15133 591 15138 647
rect 15194 591 15221 647
rect 15277 591 15303 647
rect 15359 591 15385 647
rect 15441 591 15467 647
rect 15523 591 15528 647
rect 15133 586 15528 591
rect 18585 -1026 19474 747
rect 20771 1271 21085 6537
rect 20771 1215 20776 1271
rect 20832 1215 20859 1271
rect 20915 1215 20942 1271
rect 20998 1215 21024 1271
rect 21080 1215 21085 1271
rect 20771 959 21085 1215
rect 20771 903 20776 959
rect 20832 903 20858 959
rect 20914 903 20939 959
rect 20995 903 21020 959
rect 21076 903 21085 959
rect 20771 647 21085 903
rect 20771 591 20776 647
rect 20832 591 20858 647
rect 20914 591 20939 647
rect 20995 591 21020 647
rect 21076 591 21085 647
rect 20771 503 21085 591
rect 20771 447 20776 503
rect 20832 447 20857 503
rect 20913 447 20938 503
rect 20994 447 21019 503
rect 21075 447 21085 503
rect 20771 423 21085 447
rect 20771 367 20776 423
rect 20832 367 20857 423
rect 20913 367 20938 423
rect 20994 367 21019 423
rect 21075 367 21085 423
rect 20771 362 21085 367
use sky130_fd_io__gpio_ovtv2_hotswap_guardrings  sky130_fd_io__gpio_ovtv2_hotswap_guardrings_0
timestamp 1648127584
transform 1 0 -1236 0 1 -1179
box 0 0 26980 8664
use sky130_fd_pr__pfet_01v8__example_55959141808168  sky130_fd_pr__pfet_01v8__example_55959141808168_0
timestamp 1648127584
transform 0 -1 18815 1 0 647
box -28 0 596 1489
use sky130_fd_pr__pfet_01v8__example_55959141808168  sky130_fd_pr__pfet_01v8__example_55959141808168_1
timestamp 1648127584
transform 0 -1 21965 1 0 647
box -28 0 596 1489
use sky130_fd_pr__pfet_01v8__example_55959141808168  sky130_fd_pr__pfet_01v8__example_55959141808168_2
timestamp 1648127584
transform 0 -1 15665 1 0 647
box -28 0 596 1489
use sky130_fd_pr__pfet_01v8__example_55959141808168  sky130_fd_pr__pfet_01v8__example_55959141808168_3
timestamp 1648127584
transform 0 -1 9365 1 0 647
box -28 0 596 1489
use sky130_fd_pr__pfet_01v8__example_55959141808168  sky130_fd_pr__pfet_01v8__example_55959141808168_4
timestamp 1648127584
transform 0 -1 12515 1 0 647
box -28 0 596 1489
use sky130_fd_pr__pfet_01v8__example_55959141808171  sky130_fd_pr__pfet_01v8__example_55959141808171_0
timestamp 1648127584
transform 0 -1 6215 1 0 673
box -28 0 128 1489
use sky130_fd_pr__pfet_01v8__example_55959141808171  sky130_fd_pr__pfet_01v8__example_55959141808171_1
timestamp 1648127584
transform 0 -1 3065 1 0 673
box -28 0 128 1489
use sky130_fd_pr__pfet_01v8__example_55959141808172  sky130_fd_pr__pfet_01v8__example_55959141808172_0
timestamp 1648127584
transform 0 -1 24340 1 0 1181
box -28 0 908 985
use sky130_fd_pr__pfet_01v8__example_55959141808174  sky130_fd_pr__pfet_01v8__example_55959141808174_0
timestamp 1648127584
transform 0 -1 24340 1 0 713
box -28 0 440 985
<< labels >>
flabel metal3 s 18585 1574 19474 1766 3 FreeSans 200 0 0 0 VCC_IO
port 1 nsew
flabel metal3 s 20771 1465 21085 1621 3 FreeSans 200 0 0 0 VPB_DRVR
port 2 nsew
flabel metal1 s 128 701 184 747 3 FreeSans 200 0 0 0 PSWG_H
port 3 nsew
<< properties >>
string GDS_END 39593778
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 39463704
<< end >>
