magic
tech sky130A
magscale 1 2
timestamp 1654304286
<< nwell >>
rect 30250 -2656 30362 -2335
rect 30529 -2656 30618 -2335
<< viali >>
rect 27523 -2576 27557 -2542
rect 29040 -2563 29074 -2529
rect 29208 -2563 29242 -2529
rect 29376 -2563 29410 -2529
rect 29544 -2563 29578 -2529
rect 29712 -2563 29746 -2529
rect 29880 -2563 29914 -2529
rect 30048 -2563 30082 -2529
rect 30788 -2564 30822 -2530
rect 30956 -2564 30990 -2530
rect 31124 -2564 31158 -2530
rect 31292 -2564 31326 -2530
rect 31460 -2564 31494 -2530
rect 31628 -2564 31662 -2530
rect 31796 -2564 31830 -2530
rect 27337 -2702 27371 -2668
rect 27871 -2694 27905 -2660
rect 28599 -2703 28633 -2669
rect 28800 -2698 28834 -2664
rect 28919 -2698 28953 -2664
rect 29038 -2698 29072 -2664
rect 29157 -2698 29191 -2664
rect 29276 -2698 29310 -2664
rect 29395 -2698 29429 -2664
rect 29514 -2698 29548 -2664
rect 30724 -2696 30758 -2662
rect 30843 -2696 30877 -2662
rect 30962 -2696 30996 -2662
rect 31081 -2696 31115 -2662
rect 31200 -2696 31234 -2662
rect 31319 -2696 31353 -2662
rect 31438 -2696 31472 -2662
<< metal1 >>
rect 86 1593 444 1613
rect 86 1592 386 1593
rect 86 1540 110 1592
rect 162 1541 386 1592
rect 438 1541 444 1593
rect 162 1540 444 1541
rect 86 1516 444 1540
rect 60809 851 61053 929
rect 30 -79 28869 -74
rect 30 -131 28779 -79
rect 28831 -131 28869 -79
rect 30 -135 28869 -131
rect 30628 -82 61307 -77
rect 30628 -134 30666 -82
rect 30718 -134 61307 -82
rect 30628 -138 61307 -134
rect 30 -221 26961 -216
rect 30 -273 26891 -221
rect 26943 -273 26961 -221
rect 30 -277 26961 -273
rect 32536 -224 61307 -219
rect 32536 -276 32554 -224
rect 32606 -276 61307 -224
rect 32536 -280 61307 -276
rect 30 -362 25103 -358
rect 30 -414 25004 -362
rect 25056 -414 25103 -362
rect 30 -419 25103 -414
rect 34394 -365 61307 -361
rect 34394 -417 34441 -365
rect 34493 -417 61307 -365
rect 34394 -422 61307 -417
rect 30 -503 23179 -500
rect 30 -555 23115 -503
rect 23167 -555 23179 -503
rect 30 -561 23179 -555
rect 36318 -506 61307 -503
rect 36318 -558 36330 -506
rect 36382 -558 61307 -506
rect 36318 -564 61307 -558
rect 30 -646 21303 -642
rect 30 -698 21227 -646
rect 21279 -698 21303 -646
rect 30 -703 21303 -698
rect 38194 -649 61307 -645
rect 38194 -701 38218 -649
rect 38270 -701 61307 -649
rect 38194 -706 61307 -701
rect 30 -789 19421 -784
rect 30 -841 19337 -789
rect 19389 -841 19421 -789
rect 30 -845 19421 -841
rect 40076 -792 61307 -787
rect 40076 -844 40108 -792
rect 40160 -844 61307 -792
rect 40076 -848 61307 -844
rect 30 -930 17513 -926
rect 30 -982 17451 -930
rect 17503 -982 17513 -930
rect 30 -987 17513 -982
rect 41984 -933 61307 -929
rect 41984 -985 41994 -933
rect 42046 -985 61307 -933
rect 41984 -990 61307 -985
rect 30 -1073 15637 -1068
rect 30 -1125 15563 -1073
rect 15615 -1125 15637 -1073
rect 30 -1129 15637 -1125
rect 43860 -1076 61307 -1071
rect 43860 -1128 43882 -1076
rect 43934 -1128 61307 -1076
rect 43860 -1132 61307 -1128
rect 30 -1215 13767 -1210
rect 30 -1267 13682 -1215
rect 13734 -1267 13767 -1215
rect 30 -1271 13767 -1267
rect 45730 -1218 61307 -1213
rect 45730 -1270 45763 -1218
rect 45815 -1270 61307 -1218
rect 45730 -1274 61307 -1270
rect 30 -1358 11895 -1352
rect 30 -1410 11794 -1358
rect 11846 -1410 11895 -1358
rect 30 -1413 11895 -1410
rect 47602 -1361 61307 -1355
rect 47602 -1413 47651 -1361
rect 47703 -1413 61307 -1361
rect 47602 -1416 61307 -1413
rect 30 -1500 10009 -1494
rect 30 -1552 9906 -1500
rect 9958 -1552 10009 -1500
rect 30 -1555 10009 -1552
rect 49488 -1498 59467 -1497
rect 60835 -1498 61307 -1497
rect 49488 -1503 61307 -1498
rect 49488 -1555 49539 -1503
rect 49591 -1555 61307 -1503
rect 49488 -1558 61307 -1555
rect 59370 -1559 61307 -1558
rect 30 -1642 8098 -1636
rect 30 -1694 8019 -1642
rect 8071 -1694 8098 -1642
rect 30 -1697 8098 -1694
rect 51399 -1645 61307 -1639
rect 51399 -1697 51426 -1645
rect 51478 -1697 61307 -1645
rect 51399 -1700 61307 -1697
rect 30 -1783 6222 -1778
rect 30 -1835 6129 -1783
rect 6181 -1835 6222 -1783
rect 30 -1839 6222 -1835
rect 53275 -1786 61307 -1781
rect 53275 -1838 53316 -1786
rect 53368 -1838 61307 -1786
rect 53275 -1842 61307 -1838
rect 30 -1925 4325 -1920
rect 30 -1977 4242 -1925
rect 4294 -1977 4325 -1925
rect 30 -1981 4325 -1977
rect 55172 -1928 61307 -1923
rect 55172 -1980 55203 -1928
rect 55255 -1980 61307 -1928
rect 55172 -1984 61307 -1980
rect 30 -2068 2453 -2062
rect 30 -2120 2353 -2068
rect 2405 -2120 2453 -2068
rect 30 -2123 2453 -2120
rect 57044 -2071 61307 -2065
rect 57044 -2123 57092 -2071
rect 57144 -2123 61307 -2071
rect 57044 -2126 61307 -2123
rect 30 -2209 594 -2204
rect 30 -2261 465 -2209
rect 517 -2261 594 -2209
rect 30 -2265 594 -2261
rect 58903 -2212 61307 -2207
rect 58903 -2264 58980 -2212
rect 59032 -2264 61307 -2212
rect 58903 -2268 61307 -2264
rect 30 -2351 816 -2346
rect 30 -2403 692 -2351
rect 744 -2403 816 -2351
rect 30 -2407 816 -2403
rect 27760 -2421 27836 -2325
rect 28664 -2421 28740 -2325
rect 30212 -2421 30399 -2325
rect 30491 -2421 30678 -2325
rect 59138 -2354 61307 -2349
rect 59138 -2406 59210 -2354
rect 59262 -2406 61307 -2354
rect 59138 -2410 61307 -2406
rect 30 -2490 2675 -2488
rect 30 -2542 2579 -2490
rect 2631 -2542 2675 -2490
rect 57279 -2493 61307 -2491
rect 30 -2549 2675 -2542
rect 27513 -2542 27566 -2525
rect 27513 -2576 27523 -2542
rect 27557 -2576 27566 -2542
rect 30 -2635 4586 -2630
rect 30 -2687 4468 -2635
rect 4520 -2687 4586 -2635
rect 30 -2691 4586 -2687
rect 6821 -2646 7168 -2624
rect 6821 -2658 27389 -2646
rect 6821 -2710 6910 -2658
rect 6962 -2710 7008 -2658
rect 7060 -2668 27389 -2658
rect 7060 -2702 27337 -2668
rect 27371 -2702 27389 -2668
rect 7060 -2710 27389 -2702
rect 27513 -2647 27566 -2576
rect 29028 -2529 31845 -2504
rect 29028 -2563 29040 -2529
rect 29074 -2563 29208 -2529
rect 29242 -2563 29376 -2529
rect 29410 -2563 29544 -2529
rect 29578 -2563 29712 -2529
rect 29746 -2563 29880 -2529
rect 29914 -2563 30048 -2529
rect 30082 -2530 31845 -2529
rect 30082 -2538 30788 -2530
rect 30082 -2563 30260 -2538
rect 29028 -2590 30260 -2563
rect 30312 -2590 30363 -2538
rect 30415 -2590 30466 -2538
rect 30518 -2590 30569 -2538
rect 30621 -2564 30788 -2538
rect 30822 -2564 30956 -2530
rect 30990 -2564 31124 -2530
rect 31158 -2564 31292 -2530
rect 31326 -2564 31460 -2530
rect 31494 -2564 31628 -2530
rect 31662 -2564 31796 -2530
rect 31830 -2564 31845 -2530
rect 57279 -2545 57323 -2493
rect 57375 -2545 61307 -2493
rect 57279 -2552 61307 -2545
rect 30621 -2590 31845 -2564
rect 29028 -2612 31845 -2590
rect 55368 -2638 61307 -2633
rect 27513 -2660 27923 -2647
rect 27513 -2694 27871 -2660
rect 27905 -2694 27923 -2660
rect 27513 -2708 27923 -2694
rect 28577 -2662 31768 -2653
rect 28577 -2664 30724 -2662
rect 28577 -2669 28800 -2664
rect 28577 -2703 28599 -2669
rect 28633 -2698 28800 -2669
rect 28834 -2698 28919 -2664
rect 28953 -2698 29038 -2664
rect 29072 -2698 29157 -2664
rect 29191 -2698 29276 -2664
rect 29310 -2698 29395 -2664
rect 29429 -2698 29514 -2664
rect 29548 -2696 30724 -2664
rect 30758 -2696 30843 -2662
rect 30877 -2696 30962 -2662
rect 30996 -2696 31081 -2662
rect 31115 -2696 31200 -2662
rect 31234 -2696 31319 -2662
rect 31353 -2696 31438 -2662
rect 31472 -2696 31768 -2662
rect 55368 -2690 55434 -2638
rect 55486 -2690 61307 -2638
rect 55368 -2694 61307 -2690
rect 29548 -2698 31768 -2696
rect 28633 -2703 31768 -2698
rect 28577 -2710 31768 -2703
rect 6821 -2720 27389 -2710
rect 6821 -2748 7168 -2720
rect 30 -2776 6432 -2772
rect 30 -2828 6357 -2776
rect 6409 -2828 6432 -2776
rect 30 -2833 6432 -2828
rect 53522 -2779 61307 -2775
rect 53522 -2831 53545 -2779
rect 53597 -2831 61307 -2779
rect 53522 -2836 61307 -2831
rect 30 -2920 8323 -2914
rect 30 -2972 8244 -2920
rect 8296 -2972 8323 -2920
rect 27760 -2965 27836 -2869
rect 28664 -2966 28740 -2870
rect 30212 -2965 30399 -2869
rect 30491 -2965 30678 -2869
rect 51631 -2923 61307 -2917
rect 30 -2975 8323 -2972
rect 51631 -2975 51658 -2923
rect 51710 -2975 61307 -2923
rect 51631 -2978 61307 -2975
rect 30 -3061 10211 -3056
rect 30 -3113 10132 -3061
rect 10184 -3113 10211 -3061
rect 30 -3117 10211 -3113
rect 49743 -3064 61307 -3059
rect 49743 -3116 49770 -3064
rect 49822 -3116 61307 -3064
rect 49743 -3120 61307 -3116
rect 30 -3203 12112 -3198
rect 30 -3255 12021 -3203
rect 12073 -3255 12112 -3203
rect 30 -3259 12112 -3255
rect 47842 -3206 61307 -3201
rect 47842 -3258 47881 -3206
rect 47933 -3258 61307 -3206
rect 47842 -3262 61307 -3258
rect 30 -3348 13987 -3340
rect 30 -3400 13909 -3348
rect 13961 -3400 13987 -3348
rect 30 -3401 13987 -3400
rect 45967 -3351 61307 -3343
rect 45967 -3403 45993 -3351
rect 46045 -3403 61307 -3351
rect 45967 -3404 61307 -3403
rect 30 -3487 15898 -3482
rect 30 -3539 15787 -3487
rect 15839 -3539 15898 -3487
rect 30 -3543 15898 -3539
rect 44056 -3490 61307 -3485
rect 44056 -3542 44115 -3490
rect 44167 -3542 61307 -3490
rect 44056 -3546 61307 -3542
rect 30 -3628 17796 -3624
rect 30 -3680 17678 -3628
rect 17730 -3680 17796 -3628
rect 30 -3685 17796 -3680
rect 42158 -3631 61307 -3627
rect 42158 -3683 42224 -3631
rect 42276 -3683 61307 -3631
rect 42158 -3688 61307 -3683
rect 30 -3769 19703 -3766
rect 30 -3821 19563 -3769
rect 19615 -3821 19703 -3769
rect 30 -3827 19703 -3821
rect 40251 -3772 61307 -3769
rect 40251 -3824 40339 -3772
rect 40391 -3824 61307 -3772
rect 40251 -3830 61307 -3824
rect 30 -3912 21553 -3908
rect 30 -3964 21454 -3912
rect 21506 -3964 21553 -3912
rect 30 -3969 21553 -3964
rect 38401 -3915 61307 -3911
rect 38401 -3967 38448 -3915
rect 38500 -3967 61307 -3915
rect 38401 -3972 61307 -3967
rect 30 -4055 23428 -4050
rect 30 -4107 23344 -4055
rect 23396 -4107 23428 -4055
rect 30 -4111 23428 -4107
rect 36526 -4058 61307 -4053
rect 36526 -4110 36558 -4058
rect 36610 -4110 61307 -4058
rect 36526 -4114 61307 -4110
rect 30 -4199 25325 -4192
rect 30 -4251 25227 -4199
rect 25279 -4251 25325 -4199
rect 30 -4253 25325 -4251
rect 34629 -4202 61307 -4195
rect 34629 -4254 34675 -4202
rect 34727 -4254 61307 -4202
rect 34629 -4256 61307 -4254
rect 30 -4341 27255 -4334
rect 30 -4393 27117 -4341
rect 27169 -4393 27255 -4341
rect 30 -4395 27255 -4393
rect 32699 -4344 61307 -4337
rect 32699 -4396 32785 -4344
rect 32837 -4396 61307 -4344
rect 32699 -4398 61307 -4396
rect 30 -4481 29105 -4476
rect 30 -4533 29009 -4481
rect 29061 -4533 29105 -4481
rect 30 -4537 29105 -4533
rect 30849 -4484 61307 -4479
rect 30849 -4536 30893 -4484
rect 30945 -4536 61307 -4484
rect 30849 -4540 61307 -4536
rect -167 -6186 614 -6171
rect -167 -6194 555 -6186
rect -167 -6246 -150 -6194
rect -98 -6238 555 -6194
rect 607 -6238 614 -6186
rect -98 -6246 614 -6238
rect -167 -6264 614 -6246
<< via1 >>
rect 30296 3154 30348 3206
rect 30413 3154 30465 3206
rect 30530 3154 30582 3206
rect 110 1540 162 1592
rect 386 1541 438 1593
rect 28779 -131 28831 -79
rect 30666 -134 30718 -82
rect 26891 -273 26943 -221
rect 32554 -276 32606 -224
rect 25004 -414 25056 -362
rect 34441 -417 34493 -365
rect 23115 -555 23167 -503
rect 36330 -558 36382 -506
rect 21227 -698 21279 -646
rect 38218 -701 38270 -649
rect 19337 -841 19389 -789
rect 40108 -844 40160 -792
rect 17451 -982 17503 -930
rect 41994 -985 42046 -933
rect 15563 -1125 15615 -1073
rect 43882 -1128 43934 -1076
rect 13682 -1267 13734 -1215
rect 45763 -1270 45815 -1218
rect 11794 -1410 11846 -1358
rect 47651 -1413 47703 -1361
rect 9906 -1552 9958 -1500
rect 49539 -1555 49591 -1503
rect 8019 -1694 8071 -1642
rect 51426 -1697 51478 -1645
rect 6129 -1835 6181 -1783
rect 53316 -1838 53368 -1786
rect 4242 -1977 4294 -1925
rect 55203 -1980 55255 -1928
rect 2353 -2120 2405 -2068
rect 57092 -2123 57144 -2071
rect 465 -2261 517 -2209
rect 58980 -2264 59032 -2212
rect 692 -2403 744 -2351
rect 31363 -2407 31415 -2355
rect 31493 -2407 31545 -2355
rect 31623 -2407 31675 -2355
rect 59210 -2406 59262 -2354
rect 2579 -2542 2631 -2490
rect 4468 -2687 4520 -2635
rect 6910 -2710 6962 -2658
rect 7008 -2710 7060 -2658
rect 30260 -2590 30312 -2538
rect 30363 -2590 30415 -2538
rect 30466 -2590 30518 -2538
rect 30569 -2590 30621 -2538
rect 57323 -2545 57375 -2493
rect 55434 -2690 55486 -2638
rect 6357 -2828 6409 -2776
rect 53545 -2831 53597 -2779
rect 8244 -2972 8296 -2920
rect 31353 -2937 31405 -2885
rect 31466 -2937 31518 -2885
rect 31579 -2937 31631 -2885
rect 31692 -2937 31744 -2885
rect 31805 -2937 31857 -2885
rect 51658 -2975 51710 -2923
rect 10132 -3113 10184 -3061
rect 49770 -3116 49822 -3064
rect 12021 -3255 12073 -3203
rect 47881 -3258 47933 -3206
rect 13909 -3400 13961 -3348
rect 45993 -3403 46045 -3351
rect 15787 -3539 15839 -3487
rect 44115 -3542 44167 -3490
rect 17678 -3680 17730 -3628
rect 42224 -3683 42276 -3631
rect 19563 -3821 19615 -3769
rect 40339 -3824 40391 -3772
rect 21454 -3964 21506 -3912
rect 38448 -3967 38500 -3915
rect 23344 -4107 23396 -4055
rect 36558 -4110 36610 -4058
rect 25227 -4251 25279 -4199
rect 34675 -4254 34727 -4202
rect 27117 -4393 27169 -4341
rect 32785 -4396 32837 -4344
rect 29009 -4533 29061 -4481
rect 30893 -4536 30945 -4484
rect 31353 -4826 31405 -4774
rect 31466 -4826 31518 -4774
rect 31579 -4826 31631 -4774
rect 31692 -4826 31744 -4774
rect 31805 -4826 31857 -4774
rect 31353 -4931 31405 -4879
rect 31466 -4931 31518 -4879
rect 31579 -4931 31631 -4879
rect 31692 -4931 31744 -4879
rect 31805 -4931 31857 -4879
rect -150 -6246 -98 -6194
rect 555 -6238 607 -6186
rect 30285 -9075 30337 -9023
rect 30368 -9075 30420 -9023
rect 30451 -9075 30503 -9023
rect 30534 -9075 30586 -9023
<< metal2 >>
rect 1839 6719 1883 7341
rect 3727 6719 3771 7341
rect 5615 6719 5659 7341
rect 7503 6719 7547 7341
rect 9391 6719 9435 7341
rect 11279 6719 11323 7341
rect 13167 6719 13211 7341
rect 15055 6719 15099 7341
rect 16943 6719 16987 7341
rect 18831 6719 18875 7341
rect 20719 6719 20763 7341
rect 22607 6719 22651 7341
rect 24495 6719 24539 7341
rect 26383 6719 26427 7341
rect 28271 6719 28315 7341
rect 30159 6719 30203 7341
rect 32047 6719 32091 7341
rect 33935 6719 33979 7341
rect 35823 6719 35867 7341
rect 37711 6719 37755 7341
rect 39599 6719 39643 7341
rect 41487 6719 41531 7341
rect 43375 6719 43419 7341
rect 45263 6719 45307 7341
rect 47151 6719 47195 7341
rect 49039 6719 49083 7341
rect 50927 6719 50971 7341
rect 52815 6719 52859 7341
rect 54703 6719 54747 7341
rect 56591 6719 56635 7341
rect 58479 6719 58523 7341
rect 60367 6719 60411 7341
rect 60942 6037 60978 6070
rect -159 6001 555 6037
rect 60231 6001 60978 6037
rect -159 -6171 -123 6001
rect 30232 3261 30628 3290
rect 30232 3205 30263 3261
rect 30319 3206 30372 3261
rect 30428 3206 30481 3261
rect 30537 3206 30628 3261
rect 30348 3205 30372 3206
rect 30465 3205 30481 3206
rect 30232 3159 30296 3205
rect 30348 3159 30413 3205
rect 30465 3159 30530 3205
rect 30232 3103 30263 3159
rect 30348 3154 30372 3159
rect 30465 3154 30481 3159
rect 30582 3154 30628 3206
rect 30319 3103 30372 3154
rect 30428 3103 30481 3154
rect 30537 3103 30628 3154
rect 30232 3082 30628 3103
rect 75 1592 173 1619
rect 75 1540 110 1592
rect 162 1540 173 1592
rect 75 1500 173 1540
rect 373 1593 477 1616
rect 373 1541 386 1593
rect 438 1581 477 1593
rect 60942 1581 60978 6001
rect 438 1545 649 1581
rect 60325 1545 60978 1581
rect 438 1541 477 1545
rect 373 1516 477 1541
rect -160 -6194 -49 -6171
rect -160 -6246 -150 -6194
rect -98 -6246 -49 -6194
rect -160 -6286 -49 -6246
rect 107 -10650 143 1500
rect 469 -2199 513 863
rect 2357 -2056 2401 863
rect 4245 -1916 4289 863
rect 6133 -1772 6177 863
rect 8021 -1632 8065 863
rect 9909 -1490 9953 455
rect 11797 -1348 11841 475
rect 13685 -1206 13729 465
rect 15567 -1065 15611 472
rect 17455 -924 17499 525
rect 19343 -779 19387 465
rect 21231 -636 21275 445
rect 23119 -494 23163 445
rect 25007 -353 25051 405
rect 26895 -210 26939 449
rect 28783 -64 28827 459
rect 28760 -79 28854 -64
rect 30670 -67 30714 298
rect 28760 -131 28779 -79
rect 28831 -131 28854 -79
rect 28760 -145 28854 -131
rect 30643 -82 30737 -67
rect 30643 -134 30666 -82
rect 30718 -134 30737 -82
rect 28783 -189 28827 -145
rect 30643 -148 30737 -134
rect 30670 -192 30714 -148
rect 26880 -221 26957 -210
rect 32558 -213 32602 319
rect 26880 -273 26891 -221
rect 26943 -273 26957 -221
rect 26880 -283 26957 -273
rect 32540 -224 32617 -213
rect 32540 -276 32554 -224
rect 32606 -276 32617 -224
rect 26895 -326 26939 -283
rect 32540 -286 32617 -276
rect 32558 -329 32602 -286
rect 24991 -362 25068 -353
rect 34446 -356 34490 375
rect 24991 -414 25004 -362
rect 25056 -414 25068 -362
rect 24991 -426 25068 -414
rect 34429 -365 34506 -356
rect 34429 -417 34441 -365
rect 34493 -417 34506 -365
rect 25007 -456 25051 -426
rect 34429 -429 34506 -417
rect 34446 -459 34490 -429
rect 23104 -503 23181 -494
rect 36334 -497 36378 300
rect 23104 -555 23115 -503
rect 23167 -555 23181 -503
rect 23104 -567 23181 -555
rect 36316 -506 36393 -497
rect 36316 -558 36330 -506
rect 36382 -558 36393 -506
rect 23119 -603 23163 -567
rect 36316 -570 36393 -558
rect 36334 -606 36378 -570
rect 21215 -646 21292 -636
rect 38222 -639 38266 310
rect 21215 -698 21227 -646
rect 21279 -698 21292 -646
rect 21215 -709 21292 -698
rect 38205 -649 38282 -639
rect 38205 -701 38218 -649
rect 38270 -701 38282 -649
rect 21231 -743 21275 -709
rect 38205 -712 38282 -701
rect 38222 -746 38266 -712
rect 19329 -789 19406 -779
rect 40110 -782 40154 338
rect 19329 -841 19337 -789
rect 19389 -841 19406 -789
rect 19329 -852 19406 -841
rect 40091 -792 40168 -782
rect 40091 -844 40108 -792
rect 40160 -844 40168 -792
rect 19343 -894 19387 -852
rect 40091 -855 40168 -844
rect 40110 -897 40154 -855
rect 17438 -930 17515 -924
rect 41998 -927 42042 331
rect 17438 -982 17451 -930
rect 17503 -982 17515 -930
rect 17438 -997 17515 -982
rect 41982 -933 42059 -927
rect 41982 -985 41994 -933
rect 42046 -985 42059 -933
rect 17455 -1040 17499 -997
rect 41982 -1000 42059 -985
rect 41998 -1043 42042 -1000
rect 15551 -1073 15628 -1065
rect 43886 -1068 43930 329
rect 15551 -1125 15563 -1073
rect 15615 -1125 15628 -1073
rect 15551 -1138 15628 -1125
rect 43869 -1076 43946 -1068
rect 43869 -1128 43882 -1076
rect 43934 -1128 43946 -1076
rect 15567 -1167 15611 -1138
rect 43869 -1141 43946 -1128
rect 43886 -1170 43930 -1141
rect 13670 -1215 13747 -1206
rect 45768 -1209 45812 297
rect 13670 -1267 13682 -1215
rect 13734 -1267 13747 -1215
rect 13670 -1279 13747 -1267
rect 45750 -1218 45827 -1209
rect 45750 -1270 45763 -1218
rect 45815 -1270 45827 -1218
rect 13685 -1307 13729 -1279
rect 45750 -1282 45827 -1270
rect 45768 -1310 45812 -1282
rect 11782 -1358 11859 -1348
rect 47656 -1351 47700 335
rect 11782 -1410 11794 -1358
rect 11846 -1410 11859 -1358
rect 11782 -1421 11859 -1410
rect 47638 -1361 47715 -1351
rect 47638 -1413 47651 -1361
rect 47703 -1413 47715 -1361
rect 11797 -1444 11841 -1421
rect 47638 -1424 47715 -1413
rect 47656 -1447 47700 -1424
rect 9893 -1500 9970 -1490
rect 49544 -1493 49588 320
rect 9893 -1552 9906 -1500
rect 9958 -1552 9970 -1500
rect 9893 -1563 9970 -1552
rect 49527 -1503 49604 -1493
rect 49527 -1555 49539 -1503
rect 49591 -1555 49604 -1503
rect 9909 -1601 9953 -1563
rect 49527 -1566 49604 -1555
rect 49544 -1604 49588 -1566
rect 8007 -1642 8084 -1632
rect 51432 -1635 51476 320
rect 8007 -1694 8019 -1642
rect 8071 -1694 8084 -1642
rect 8007 -1705 8084 -1694
rect 51413 -1645 51490 -1635
rect 51413 -1697 51426 -1645
rect 51478 -1697 51490 -1645
rect 8021 -1738 8065 -1705
rect 51413 -1708 51490 -1697
rect 51432 -1741 51476 -1708
rect 6119 -1783 6196 -1772
rect 53320 -1775 53364 333
rect 6119 -1835 6129 -1783
rect 6181 -1835 6196 -1783
rect 6119 -1845 6196 -1835
rect 53301 -1786 53378 -1775
rect 53301 -1838 53316 -1786
rect 53368 -1838 53378 -1786
rect 6133 -1881 6177 -1845
rect 53301 -1848 53378 -1838
rect 4229 -1925 4306 -1916
rect 4229 -1977 4242 -1925
rect 4294 -1977 4306 -1925
rect 4229 -1989 4306 -1977
rect 30233 -1921 30630 -1882
rect 53320 -1884 53364 -1848
rect 55208 -1919 55252 350
rect 30233 -1977 30256 -1921
rect 30312 -1977 30360 -1921
rect 30416 -1977 30464 -1921
rect 30520 -1977 30568 -1921
rect 30624 -1977 30630 -1921
rect 4245 -2028 4289 -1989
rect 30233 -2020 30630 -1977
rect 55191 -1928 55268 -1919
rect 55191 -1980 55203 -1928
rect 55255 -1980 55268 -1928
rect 55191 -1992 55268 -1980
rect 2345 -2068 2422 -2056
rect 2345 -2120 2353 -2068
rect 2405 -2120 2422 -2068
rect 2345 -2129 2422 -2120
rect 30233 -2076 30256 -2020
rect 30312 -2076 30360 -2020
rect 30416 -2076 30464 -2020
rect 30520 -2076 30568 -2020
rect 30624 -2076 30630 -2020
rect 55208 -2031 55252 -1992
rect 57096 -2059 57140 348
rect 2357 -2165 2401 -2129
rect 452 -2209 529 -2199
rect 452 -2261 465 -2209
rect 517 -2261 529 -2209
rect 452 -2272 529 -2261
rect 469 -2295 513 -2272
rect 698 -2340 742 -2310
rect 681 -2351 760 -2340
rect 681 -2403 692 -2351
rect 744 -2403 760 -2351
rect 681 -2416 760 -2403
rect 698 -5048 742 -2416
rect 2586 -2481 2630 -2437
rect 2567 -2490 2646 -2481
rect 2567 -2542 2579 -2490
rect 2631 -2542 2646 -2490
rect 2567 -2557 2646 -2542
rect 30233 -2538 30630 -2076
rect 57075 -2071 57152 -2059
rect 57075 -2123 57092 -2071
rect 57144 -2123 57152 -2071
rect 57075 -2132 57152 -2123
rect 57096 -2168 57140 -2132
rect 58984 -2202 59028 346
rect 58968 -2212 59045 -2202
rect 58968 -2264 58980 -2212
rect 59032 -2264 59045 -2212
rect 58968 -2275 59045 -2264
rect 58984 -2298 59028 -2275
rect 31324 -2351 31725 -2326
rect 59212 -2343 59256 -2313
rect 31324 -2407 31363 -2351
rect 31419 -2407 31492 -2351
rect 31548 -2407 31621 -2351
rect 31677 -2407 31725 -2351
rect 31324 -2420 31725 -2407
rect 59194 -2354 59273 -2343
rect 59194 -2406 59210 -2354
rect 59262 -2406 59273 -2354
rect 59194 -2419 59273 -2406
rect 57324 -2484 57368 -2440
rect 2586 -5094 2630 -2557
rect 4474 -2627 4518 -2554
rect 30233 -2590 30260 -2538
rect 30312 -2590 30363 -2538
rect 30415 -2590 30466 -2538
rect 30518 -2590 30569 -2538
rect 30621 -2590 30630 -2538
rect 57308 -2493 57387 -2484
rect 57308 -2545 57323 -2493
rect 57375 -2545 57387 -2493
rect 4449 -2635 4528 -2627
rect 4449 -2687 4468 -2635
rect 4520 -2687 4528 -2635
rect 4449 -2703 4528 -2687
rect 6821 -2654 7168 -2624
rect 6821 -2658 6911 -2654
rect 4474 -5131 4518 -2703
rect 6362 -2768 6406 -2694
rect 6821 -2710 6910 -2658
rect 6967 -2710 7008 -2654
rect 7064 -2710 7168 -2654
rect 6821 -2748 7168 -2710
rect 6344 -2776 6423 -2768
rect 6344 -2828 6357 -2776
rect 6409 -2828 6423 -2776
rect 6344 -2844 6423 -2828
rect 6362 -5082 6406 -2844
rect 8250 -2909 8294 -2860
rect 8233 -2920 8312 -2909
rect 8233 -2972 8244 -2920
rect 8296 -2972 8312 -2920
rect 8233 -2985 8312 -2972
rect 8250 -5045 8294 -2985
rect 10138 -3051 10182 -3006
rect 10121 -3061 10200 -3051
rect 10121 -3113 10132 -3061
rect 10184 -3113 10200 -3061
rect 10121 -3127 10200 -3113
rect 10138 -5082 10182 -3127
rect 12026 -3194 12070 -3153
rect 12010 -3203 12089 -3194
rect 12010 -3255 12021 -3203
rect 12073 -3255 12089 -3203
rect 12010 -3270 12089 -3255
rect 30233 -3250 30630 -2590
rect 55436 -2630 55480 -2557
rect 57308 -2560 57387 -2545
rect 55426 -2638 55505 -2630
rect 55426 -2690 55434 -2638
rect 55486 -2690 55505 -2638
rect 53548 -2771 53592 -2697
rect 55426 -2706 55505 -2690
rect 53531 -2779 53610 -2771
rect 53531 -2831 53545 -2779
rect 53597 -2831 53610 -2779
rect 53531 -2847 53610 -2831
rect 12026 -5106 12070 -3270
rect 30233 -3306 30269 -3250
rect 30325 -3306 30357 -3250
rect 30413 -3306 30445 -3250
rect 30501 -3306 30533 -3250
rect 30589 -3306 30630 -3250
rect 13914 -3339 13958 -3312
rect 13898 -3348 13977 -3339
rect 13898 -3400 13909 -3348
rect 13961 -3400 13977 -3348
rect 13898 -3415 13977 -3400
rect 30233 -3345 30630 -3306
rect 30233 -3401 30269 -3345
rect 30325 -3401 30357 -3345
rect 30413 -3401 30445 -3345
rect 30501 -3401 30533 -3345
rect 30589 -3401 30630 -3345
rect 13914 -5082 13958 -3415
rect 30233 -3432 30630 -3401
rect 31298 -2885 31965 -2868
rect 31298 -2937 31353 -2885
rect 31405 -2937 31466 -2885
rect 31518 -2937 31579 -2885
rect 31631 -2937 31692 -2885
rect 31744 -2937 31805 -2885
rect 31857 -2937 31965 -2885
rect 51660 -2912 51704 -2863
rect 15796 -3477 15840 -3435
rect 15776 -3487 15855 -3477
rect 15776 -3539 15787 -3487
rect 15839 -3539 15855 -3487
rect 15776 -3553 15855 -3539
rect 15796 -5137 15840 -3553
rect 17684 -3619 17728 -3563
rect 17666 -3628 17745 -3619
rect 17666 -3680 17678 -3628
rect 17730 -3680 17745 -3628
rect 17666 -3695 17745 -3680
rect 17684 -5106 17728 -3695
rect 19572 -3760 19616 -3704
rect 19552 -3769 19631 -3760
rect 19552 -3821 19563 -3769
rect 19615 -3821 19631 -3769
rect 19552 -3836 19631 -3821
rect 19572 -5064 19616 -3836
rect 21460 -3902 21504 -3845
rect 21442 -3912 21521 -3902
rect 21442 -3964 21454 -3912
rect 21506 -3964 21521 -3912
rect 21442 -3978 21521 -3964
rect 21460 -5088 21504 -3978
rect 23348 -4045 23392 -3979
rect 23332 -4055 23411 -4045
rect 23332 -4107 23344 -4055
rect 23396 -4107 23411 -4055
rect 23332 -4121 23411 -4107
rect 23348 -5137 23392 -4121
rect 25236 -4186 25280 -4132
rect 25214 -4199 25293 -4186
rect 25214 -4251 25227 -4199
rect 25279 -4251 25293 -4199
rect 25214 -4262 25293 -4251
rect 25236 -5106 25280 -4262
rect 27124 -4328 27168 -4291
rect 27108 -4341 27187 -4328
rect 27108 -4393 27117 -4341
rect 27169 -4393 27187 -4341
rect 27108 -4404 27187 -4393
rect 27124 -5106 27168 -4404
rect 29012 -4470 29056 -4395
rect 28998 -4481 29077 -4470
rect 30898 -4473 30942 -4398
rect 28998 -4533 29009 -4481
rect 29061 -4533 29077 -4481
rect 28998 -4546 29077 -4533
rect 30877 -4484 30956 -4473
rect 30877 -4536 30893 -4484
rect 30945 -4536 30956 -4484
rect 29012 -5100 29056 -4546
rect 30877 -4549 30956 -4536
rect 30898 -5005 30942 -4549
rect 31298 -4774 31965 -2937
rect 51642 -2923 51721 -2912
rect 51642 -2975 51658 -2923
rect 51710 -2975 51721 -2923
rect 51642 -2988 51721 -2975
rect 49772 -3054 49816 -3009
rect 49754 -3064 49833 -3054
rect 49754 -3116 49770 -3064
rect 49822 -3116 49833 -3064
rect 49754 -3130 49833 -3116
rect 47884 -3197 47928 -3156
rect 47865 -3206 47944 -3197
rect 47865 -3258 47881 -3206
rect 47933 -3258 47944 -3206
rect 47865 -3273 47944 -3258
rect 45996 -3342 46040 -3315
rect 45977 -3351 46056 -3342
rect 45977 -3403 45993 -3351
rect 46045 -3403 46056 -3351
rect 45977 -3418 46056 -3403
rect 44114 -3480 44158 -3438
rect 44099 -3490 44178 -3480
rect 44099 -3542 44115 -3490
rect 44167 -3542 44178 -3490
rect 44099 -3556 44178 -3542
rect 42226 -3622 42270 -3566
rect 42209 -3631 42288 -3622
rect 42209 -3683 42224 -3631
rect 42276 -3683 42288 -3631
rect 42209 -3698 42288 -3683
rect 40338 -3763 40382 -3707
rect 40323 -3772 40402 -3763
rect 40323 -3824 40339 -3772
rect 40391 -3824 40402 -3772
rect 40323 -3839 40402 -3824
rect 38450 -3905 38494 -3848
rect 38433 -3915 38512 -3905
rect 38433 -3967 38448 -3915
rect 38500 -3967 38512 -3915
rect 38433 -3981 38512 -3967
rect 36562 -4048 36606 -3982
rect 36543 -4058 36622 -4048
rect 36543 -4110 36558 -4058
rect 36610 -4110 36622 -4058
rect 36543 -4124 36622 -4110
rect 34674 -4189 34718 -4135
rect 34661 -4202 34740 -4189
rect 34661 -4254 34675 -4202
rect 34727 -4254 34740 -4202
rect 34661 -4265 34740 -4254
rect 32786 -4331 32830 -4294
rect 32767 -4344 32846 -4331
rect 32767 -4396 32785 -4344
rect 32837 -4396 32846 -4344
rect 32767 -4407 32846 -4396
rect 31298 -4826 31353 -4774
rect 31405 -4826 31466 -4774
rect 31518 -4826 31579 -4774
rect 31631 -4826 31692 -4774
rect 31744 -4826 31805 -4774
rect 31857 -4826 31965 -4774
rect 31298 -4879 31965 -4826
rect 31298 -4931 31353 -4879
rect 31405 -4931 31466 -4879
rect 31518 -4931 31579 -4879
rect 31631 -4931 31692 -4879
rect 31744 -4931 31805 -4879
rect 31857 -4931 31965 -4879
rect 31298 -4979 31965 -4931
rect 32786 -4958 32830 -4407
rect 34674 -4996 34718 -4265
rect 36562 -4999 36606 -4124
rect 38450 -5005 38494 -3981
rect 40338 -4979 40382 -3839
rect 42226 -5054 42270 -3698
rect 44114 -5011 44158 -3556
rect 45996 -4992 46040 -3418
rect 47884 -5028 47928 -3273
rect 49772 -5039 49816 -3130
rect 51660 -5013 51704 -2988
rect 53548 -4988 53592 -2847
rect 55436 -5030 55480 -2706
rect 57324 -4969 57368 -2560
rect 59212 -4999 59256 -2419
rect 548 -6186 618 -6165
rect 548 -6238 555 -6186
rect 607 -6194 618 -6186
rect 607 -6230 878 -6194
rect 60554 -6230 61279 -6194
rect 607 -6238 618 -6230
rect 548 -6269 618 -6238
rect 30233 -8974 30630 -8941
rect 30233 -9030 30274 -8974
rect 30330 -9023 30366 -8974
rect 30422 -9023 30458 -8974
rect 30514 -9023 30550 -8974
rect 30337 -9030 30366 -9023
rect 30422 -9030 30451 -9023
rect 30514 -9030 30534 -9023
rect 30606 -9030 30630 -8974
rect 30233 -9065 30285 -9030
rect 30337 -9065 30368 -9030
rect 30420 -9065 30451 -9030
rect 30503 -9065 30534 -9030
rect 30586 -9065 30630 -9030
rect 30233 -9121 30274 -9065
rect 30337 -9075 30366 -9065
rect 30422 -9075 30451 -9065
rect 30514 -9075 30534 -9065
rect 30330 -9121 30366 -9075
rect 30422 -9121 30458 -9075
rect 30514 -9121 30550 -9075
rect 30606 -9121 30630 -9065
rect 30233 -9147 30630 -9121
rect 61243 -10650 61279 -6230
rect 107 -10686 784 -10650
rect 60460 -10686 61279 -10650
rect 61243 -10697 61279 -10686
rect 2068 -11990 2112 -11368
rect 3956 -11990 4000 -11368
rect 5844 -11990 5888 -11368
rect 7732 -11990 7776 -11368
rect 9620 -11990 9664 -11368
rect 11508 -11990 11552 -11368
rect 13396 -11990 13440 -11368
rect 15284 -11990 15328 -11368
rect 17172 -11990 17216 -11368
rect 19060 -11990 19104 -11368
rect 20948 -11990 20992 -11368
rect 22836 -11990 22880 -11368
rect 24724 -11990 24768 -11368
rect 26612 -11990 26656 -11368
rect 28500 -11990 28544 -11368
rect 30388 -11990 30432 -11368
rect 32276 -11990 32320 -11368
rect 34164 -11990 34208 -11368
rect 36052 -11990 36096 -11368
rect 37940 -11990 37984 -11368
rect 39828 -11990 39872 -11368
rect 41716 -11990 41760 -11368
rect 43604 -11990 43648 -11368
rect 45492 -11990 45536 -11368
rect 47380 -11990 47424 -11368
rect 49268 -11990 49312 -11368
rect 51156 -11990 51200 -11368
rect 53044 -11990 53088 -11368
rect 54932 -11990 54976 -11368
rect 56820 -11990 56864 -11368
rect 58708 -11990 58752 -11368
rect 60596 -11990 60640 -11368
<< via2 >>
rect 30263 3206 30319 3261
rect 30372 3206 30428 3261
rect 30481 3206 30537 3261
rect 30263 3205 30296 3206
rect 30296 3205 30319 3206
rect 30372 3205 30413 3206
rect 30413 3205 30428 3206
rect 30481 3205 30530 3206
rect 30530 3205 30537 3206
rect 30263 3154 30296 3159
rect 30296 3154 30319 3159
rect 30372 3154 30413 3159
rect 30413 3154 30428 3159
rect 30481 3154 30530 3159
rect 30530 3154 30537 3159
rect 30263 3103 30319 3154
rect 30372 3103 30428 3154
rect 30481 3103 30537 3154
rect 30256 -1977 30312 -1921
rect 30360 -1977 30416 -1921
rect 30464 -1977 30520 -1921
rect 30568 -1977 30624 -1921
rect 30256 -2076 30312 -2020
rect 30360 -2076 30416 -2020
rect 30464 -2076 30520 -2020
rect 30568 -2076 30624 -2020
rect 31363 -2355 31419 -2351
rect 31363 -2407 31415 -2355
rect 31415 -2407 31419 -2355
rect 31492 -2355 31548 -2351
rect 31492 -2407 31493 -2355
rect 31493 -2407 31545 -2355
rect 31545 -2407 31548 -2355
rect 31621 -2355 31677 -2351
rect 31621 -2407 31623 -2355
rect 31623 -2407 31675 -2355
rect 31675 -2407 31677 -2355
rect 6911 -2658 6967 -2654
rect 6911 -2710 6962 -2658
rect 6962 -2710 6967 -2658
rect 7008 -2658 7064 -2654
rect 7008 -2710 7060 -2658
rect 7060 -2710 7064 -2658
rect 30269 -3306 30325 -3250
rect 30357 -3306 30413 -3250
rect 30445 -3306 30501 -3250
rect 30533 -3306 30589 -3250
rect 30269 -3401 30325 -3345
rect 30357 -3401 30413 -3345
rect 30445 -3401 30501 -3345
rect 30533 -3401 30589 -3345
rect 30274 -9023 30330 -8974
rect 30366 -9023 30422 -8974
rect 30458 -9023 30514 -8974
rect 30550 -9023 30606 -8974
rect 30274 -9030 30285 -9023
rect 30285 -9030 30330 -9023
rect 30366 -9030 30368 -9023
rect 30368 -9030 30420 -9023
rect 30420 -9030 30422 -9023
rect 30458 -9030 30503 -9023
rect 30503 -9030 30514 -9023
rect 30550 -9030 30586 -9023
rect 30586 -9030 30606 -9023
rect 30274 -9075 30285 -9065
rect 30285 -9075 30330 -9065
rect 30366 -9075 30368 -9065
rect 30368 -9075 30420 -9065
rect 30420 -9075 30422 -9065
rect 30458 -9075 30503 -9065
rect 30503 -9075 30514 -9065
rect 30550 -9075 30586 -9065
rect 30586 -9075 30606 -9065
rect 30274 -9121 30330 -9075
rect 30366 -9121 30422 -9075
rect 30458 -9121 30514 -9075
rect 30550 -9121 30606 -9075
<< metal3 >>
rect 30232 3261 30627 3290
rect 30232 3205 30263 3261
rect 30319 3238 30372 3261
rect 30428 3205 30481 3261
rect 30537 3205 30627 3261
rect 30232 3159 30306 3205
rect 30402 3159 30627 3205
rect 30232 3103 30263 3159
rect 30319 3103 30372 3130
rect 30428 3103 30481 3159
rect 30537 3103 30627 3159
rect 30232 3082 30627 3103
rect 30232 -1921 30629 -1879
rect 30232 -1977 30256 -1921
rect 30312 -1946 30360 -1921
rect 30416 -1977 30464 -1921
rect 30520 -1946 30568 -1921
rect 30624 -1977 30629 -1921
rect 30232 -2020 30297 -1977
rect 30393 -2020 30479 -1977
rect 30575 -2020 30629 -1977
rect 30232 -2076 30256 -2020
rect 30312 -2076 30360 -2054
rect 30416 -2076 30464 -2020
rect 30520 -2076 30568 -2054
rect 30624 -2076 30629 -2020
rect 30232 -2103 30629 -2076
rect 31324 -2337 31725 -2326
rect 31324 -2351 31445 -2337
rect 31619 -2351 31725 -2337
rect 31324 -2407 31363 -2351
rect 31419 -2401 31445 -2351
rect 31619 -2401 31621 -2351
rect 31419 -2407 31492 -2401
rect 31548 -2407 31621 -2401
rect 31677 -2407 31725 -2351
rect 31324 -2420 31725 -2407
rect 6821 -2638 7168 -2624
rect -280 -2654 7168 -2638
rect -280 -2710 6911 -2654
rect 6967 -2710 7008 -2654
rect 7064 -2710 7168 -2654
rect -280 -2728 7168 -2710
rect 6821 -2748 7168 -2728
rect 30233 -3250 30630 -3192
rect 30233 -3306 30269 -3250
rect 30325 -3269 30357 -3250
rect 30413 -3306 30445 -3250
rect 30501 -3269 30533 -3250
rect 30589 -3306 30630 -3250
rect 30233 -3345 30289 -3306
rect 30385 -3345 30479 -3306
rect 30575 -3345 30630 -3306
rect 30233 -3401 30269 -3345
rect 30325 -3401 30357 -3377
rect 30413 -3401 30445 -3345
rect 30501 -3401 30533 -3377
rect 30589 -3401 30630 -3345
rect 30233 -3432 30630 -3401
rect 30233 -8974 30630 -8941
rect 30233 -9030 30274 -8974
rect 30330 -8998 30366 -8974
rect 30422 -9030 30458 -8974
rect 30514 -8997 30550 -8974
rect 30606 -9030 30630 -8974
rect 30233 -9065 30301 -9030
rect 30397 -9065 30475 -9030
rect 30571 -9065 30630 -9030
rect 30233 -9121 30274 -9065
rect 30330 -9121 30366 -9106
rect 30422 -9121 30458 -9065
rect 30514 -9121 30550 -9105
rect 30606 -9121 30630 -9065
rect 30233 -9147 30630 -9121
<< via3 >>
rect 30306 3205 30319 3238
rect 30319 3205 30372 3238
rect 30372 3205 30402 3238
rect 30306 3159 30402 3205
rect 30306 3130 30319 3159
rect 30319 3130 30372 3159
rect 30372 3130 30402 3159
rect 31369 2236 31493 2402
rect 31568 2236 31692 2402
rect 30297 -1977 30312 -1946
rect 30312 -1977 30360 -1946
rect 30360 -1977 30393 -1946
rect 30479 -1977 30520 -1946
rect 30520 -1977 30568 -1946
rect 30568 -1977 30575 -1946
rect 30297 -2020 30393 -1977
rect 30479 -2020 30575 -1977
rect 30297 -2054 30312 -2020
rect 30312 -2054 30360 -2020
rect 30360 -2054 30393 -2020
rect 30479 -2054 30520 -2020
rect 30520 -2054 30568 -2020
rect 30568 -2054 30575 -2020
rect 31445 -2351 31619 -2337
rect 31445 -2401 31492 -2351
rect 31492 -2401 31548 -2351
rect 31548 -2401 31619 -2351
rect 30289 -3306 30325 -3269
rect 30325 -3306 30357 -3269
rect 30357 -3306 30385 -3269
rect 30479 -3306 30501 -3269
rect 30501 -3306 30533 -3269
rect 30533 -3306 30575 -3269
rect 30289 -3345 30385 -3306
rect 30479 -3345 30575 -3306
rect 30289 -3377 30325 -3345
rect 30325 -3377 30357 -3345
rect 30357 -3377 30385 -3345
rect 30479 -3377 30501 -3345
rect 30501 -3377 30533 -3345
rect 30533 -3377 30575 -3345
rect 2976 -4948 3082 -4770
rect 3178 -4948 3284 -4770
rect 3364 -4948 3470 -4770
rect 3544 -4948 3650 -4770
rect 1754 -7084 1860 -6906
rect 1932 -7084 2038 -6906
rect 2108 -7084 2214 -6906
rect 30301 -9030 30330 -8998
rect 30330 -9030 30366 -8998
rect 30366 -9030 30397 -8998
rect 30475 -9030 30514 -8997
rect 30514 -9030 30550 -8997
rect 30550 -9030 30571 -8997
rect 30301 -9065 30397 -9030
rect 30475 -9065 30571 -9030
rect 30301 -9106 30330 -9065
rect 30330 -9106 30366 -9065
rect 30366 -9106 30397 -9065
rect 30475 -9105 30514 -9065
rect 30514 -9105 30550 -9065
rect 30550 -9105 30571 -9065
rect 1758 -10020 1864 -9842
rect 1918 -10020 2024 -9842
rect 2078 -10022 2184 -9844
rect 3012 -12122 3118 -11944
rect 3210 -12122 3316 -11944
rect 3410 -12122 3516 -11944
<< metal4 >>
rect 1683 -6906 2301 5164
rect 1683 -7084 1754 -6906
rect 1860 -7084 1932 -6906
rect 2038 -7084 2108 -6906
rect 2214 -7084 2301 -6906
rect 1683 -9842 2301 -7084
rect 1683 -10020 1758 -9842
rect 1864 -10020 1918 -9842
rect 2024 -9844 2301 -9842
rect 2024 -10020 2078 -9844
rect 1683 -10022 2078 -10020
rect 2184 -10022 2301 -9844
rect 1683 -10223 2301 -10022
rect 2916 -4770 3700 3798
rect 30232 3238 30629 3350
rect 30232 3130 30306 3238
rect 30402 3130 30629 3238
rect 30232 -1442 30629 3130
rect 30231 -1803 30629 -1442
rect 30232 -1946 30629 -1803
rect 30232 -2054 30297 -1946
rect 30393 -2054 30479 -1946
rect 30575 -2054 30629 -1946
rect 30232 -2103 30629 -2054
rect 31317 2402 31721 2521
rect 31317 2236 31369 2402
rect 31493 2236 31568 2402
rect 31692 2236 31721 2402
rect 31317 -2309 31721 2236
rect 31317 -2331 31725 -2309
rect 31324 -2337 31725 -2331
rect 31324 -2401 31445 -2337
rect 31619 -2401 31725 -2337
rect 31324 -2420 31725 -2401
rect 2916 -4948 2976 -4770
rect 3082 -4948 3178 -4770
rect 3284 -4948 3364 -4770
rect 3470 -4948 3544 -4770
rect 3650 -4948 3700 -4770
rect 2916 -11944 3700 -4948
rect 30234 -3269 30630 -3193
rect 30234 -3377 30289 -3269
rect 30385 -3377 30479 -3269
rect 30575 -3377 30630 -3269
rect 30234 -8997 30630 -3377
rect 30234 -8998 30475 -8997
rect 30234 -9106 30301 -8998
rect 30397 -9105 30475 -8998
rect 30571 -9105 30630 -8997
rect 30397 -9106 30630 -9105
rect 30234 -9209 30630 -9106
rect 2916 -12122 3012 -11944
rect 3118 -12122 3210 -11944
rect 3316 -12122 3410 -11944
rect 3516 -12122 3700 -11944
rect 2916 -12224 3700 -12122
use BR128half  BR128half_0
timestamp 1654224521
transform 1 0 449 0 1 71
box -430 -58 60604 7443
use BR128half  BR128half_1
timestamp 1654224521
transform -1 0 60660 0 1 -12160
box -430 -58 60604 7443
use sky130_fd_sc_hd__buf_2  sky130_fd_sc_hd__buf_2_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 27300 0 1 -2917
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0
timestamp 1650294714
transform 1 0 27836 0 1 -2917
box -38 -48 866 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0 ~/open-puf/layout
timestamp 1654066915
transform 1 0 28740 0 1 -2917
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_1
timestamp 1654066915
transform 1 0 30656 0 1 -2917
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDK_ROOT/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1650294714
transform 1 0 30399 0 1 -2917
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1650294714
transform 1 0 27668 0 1 -2917
box -38 -48 130 592
<< labels >>
flabel metal4 1683 -6906 2301 5164 1 FreeSans 1600 0 0 0 VDD
flabel space 2916 -4770 3700 7281 1 FreeSans 1600 0 0 0 VSS
flabel metal1 60809 851 61053 929 1 FreeSans 800 0 0 0 OUT
flabel metal2 60367 6719 60411 7341 1 FreeSans 1200 0 0 0 C[0]
flabel metal2 58479 6719 58523 7341 1 FreeSans 1200 0 0 0 C[1]
flabel metal2 56591 6719 56635 7341 1 FreeSans 1200 0 0 0 C[2]
flabel metal2 54703 6719 54747 7341 1 FreeSans 1200 0 0 0 C[3]
flabel metal2 52815 6719 52859 7341 1 FreeSans 1200 0 0 0 C[4]
flabel metal2 50927 6719 50971 7341 1 FreeSans 1200 0 0 0 C[5]
flabel metal2 49039 6719 49083 7341 1 FreeSans 1200 0 0 0 C[6]
flabel metal2 47151 6719 47195 7341 1 FreeSans 1200 0 0 0 C[7]
flabel metal2 45263 6719 45307 7341 1 FreeSans 1200 0 0 0 C[8]
flabel metal2 43375 6719 43419 7341 1 FreeSans 1200 0 0 0 C[9]
flabel metal2 41487 6719 41531 7341 1 FreeSans 1200 0 0 0 C[10]
flabel metal2 39599 6719 39643 7341 1 FreeSans 1200 0 0 0 C[11]
flabel metal2 37711 6719 37755 7341 1 FreeSans 1200 0 0 0 C[12]
flabel metal2 35823 6719 35867 7341 1 FreeSans 1200 0 0 0 C[13]
flabel metal2 33935 6719 33979 7341 1 FreeSans 1200 0 0 0 C[14]
flabel metal2 32047 6719 32091 7341 1 FreeSans 1200 0 0 0 C[15]
flabel metal2 30159 6719 30203 7341 1 FreeSans 1200 0 0 0 C[16]
flabel metal2 28271 6719 28315 7341 1 FreeSans 1200 0 0 0 C[17]
flabel metal2 26383 6719 26427 7341 1 FreeSans 1200 0 0 0 C[18]
flabel metal2 24495 6719 24539 7341 1 FreeSans 1200 0 0 0 C[19]
flabel metal2 22607 6719 22651 7341 1 FreeSans 1200 0 0 0 C[20]
flabel metal2 20719 6719 20763 7341 1 FreeSans 1200 0 0 0 C[21]
flabel metal2 18831 6719 18875 7341 1 FreeSans 1200 0 0 0 C[22]
flabel metal2 16943 6719 16987 7341 1 FreeSans 1200 0 0 0 C[23]
flabel metal2 15055 6719 15099 7341 1 FreeSans 1200 0 0 0 C[24]
flabel metal2 13167 6719 13211 7341 1 FreeSans 1200 0 0 0 C[25]
flabel metal2 11279 6719 11323 7341 1 FreeSans 1200 0 0 0 C[26]
flabel metal2 9391 6719 9435 7341 1 FreeSans 1200 0 0 0 C[27]
flabel metal2 7503 6719 7547 7341 1 FreeSans 1200 0 0 0 C[28]
flabel metal2 5615 6719 5659 7341 1 FreeSans 1200 0 0 0 C[29]
flabel metal2 3727 6719 3771 7341 1 FreeSans 1200 0 0 0 C[30]
flabel metal2 1839 6719 1883 7341 1 FreeSans 1200 0 0 0 C[31]
flabel metal2 60596 -11990 60640 -11368 1 FreeSans 1200 0 0 0 C[64]
flabel metal2 58708 -11990 58752 -11368 1 FreeSans 1200 0 0 0 C[65]
flabel metal2 56820 -11990 56864 -11368 1 FreeSans 1200 0 0 0 C[66]
flabel metal2 54932 -11990 54976 -11368 1 FreeSans 1200 0 0 0 C[67]
flabel metal2 53044 -11990 53088 -11368 1 FreeSans 1200 0 0 0 C[68]
flabel metal2 51156 -11990 51200 -11368 1 FreeSans 1200 0 0 0 C[69]
flabel metal2 49268 -11990 49312 -11368 1 FreeSans 1200 0 0 0 C[70]
flabel metal2 47380 -11990 47424 -11368 1 FreeSans 1200 0 0 0 C[71]
flabel metal2 45492 -11990 45536 -11368 1 FreeSans 1200 0 0 0 C[72]
flabel metal2 43604 -11990 43648 -11368 1 FreeSans 1200 0 0 0 C[73]
flabel metal2 41716 -11990 41760 -11368 1 FreeSans 1200 0 0 0 C[74]
flabel metal2 39828 -11990 39872 -11368 1 FreeSans 1200 0 0 0 C[75]
flabel metal2 37940 -11990 37984 -11368 1 FreeSans 1200 0 0 0 C[76]
flabel metal2 36052 -11990 36096 -11368 1 FreeSans 1200 0 0 0 C[77]
flabel metal2 34164 -11990 34208 -11368 1 FreeSans 1200 0 0 0 C[78]
flabel metal2 32276 -11990 32320 -11368 1 FreeSans 1200 0 0 0 C[79]
flabel metal2 30388 -11990 30432 -11368 1 FreeSans 1200 0 0 0 C[80]
flabel metal2 28500 -11990 28544 -11368 1 FreeSans 1200 0 0 0 C[81]
flabel metal2 26612 -11990 26656 -11368 1 FreeSans 1200 0 0 0 C[82]
flabel metal2 24724 -11990 24768 -11368 1 FreeSans 1200 0 0 0 C[83]
flabel metal2 22836 -11990 22880 -11368 1 FreeSans 1200 0 0 0 C[84]
flabel metal2 20948 -11990 20992 -11368 1 FreeSans 1200 0 0 0 C[85]
flabel metal2 19060 -11990 19104 -11368 1 FreeSans 1200 0 0 0 C[86]
flabel metal2 17172 -11990 17216 -11368 1 FreeSans 1200 0 0 0 C[87]
flabel metal2 15284 -11990 15328 -11368 1 FreeSans 1200 0 0 0 C[88]
flabel metal2 13396 -11990 13440 -11368 1 FreeSans 1200 0 0 0 C[89]
flabel metal2 11508 -11990 11552 -11368 1 FreeSans 1200 0 0 0 C[90]
flabel metal2 9620 -11990 9664 -11368 1 FreeSans 1200 0 0 0 C[91]
flabel metal2 7732 -11990 7776 -11368 1 FreeSans 1200 0 0 0 C[92]
flabel metal2 5844 -11990 5888 -11368 1 FreeSans 1200 0 0 0 C[93]
flabel metal2 3956 -11990 4000 -11368 1 FreeSans 1200 0 0 0 C[94]
flabel metal2 2068 -11990 2112 -11368 1 FreeSans 1200 0 0 0 C[95]
flabel metal1 30 -135 438 -74 1 FreeSans 800 0 0 0 C[111]
flabel metal1 30 -277 438 -216 1 FreeSans 800 0 0 0 C[110]
flabel metal1 30 -419 438 -358 1 FreeSans 800 0 0 0 C[109]
flabel metal1 30 -561 438 -500 1 FreeSans 800 0 0 0 C[108]
flabel metal1 30 -703 438 -642 1 FreeSans 800 0 0 0 C[107]
flabel metal1 30 -845 438 -784 1 FreeSans 800 0 0 0 C[106]
flabel metal1 30 -987 438 -926 1 FreeSans 800 0 0 0 C[105]
flabel metal1 30 -1129 438 -1068 1 FreeSans 800 0 0 0 C[104]
flabel metal1 30 -1271 438 -1210 1 FreeSans 800 0 0 0 C[103]
flabel metal1 30 -1413 438 -1352 1 FreeSans 800 0 0 0 C[102]
flabel metal1 30 -1555 438 -1494 1 FreeSans 800 0 0 0 C[101]
flabel metal1 30 -1697 438 -1636 1 FreeSans 800 0 0 0 C[100]
flabel metal1 30 -1839 438 -1778 1 FreeSans 800 0 0 0 C[99]
flabel metal1 30 -1981 438 -1920 1 FreeSans 800 0 0 0 C[98]
flabel metal1 30 -2123 438 -2062 1 FreeSans 800 0 0 0 C[97]
flabel metal1 30 -2265 438 -2204 1 FreeSans 800 0 0 0 C[96]
flabel metal1 30 -2407 438 -2346 1 FreeSans 800 0 0 0 C[32]
flabel metal1 30 -2549 438 -2488 1 FreeSans 800 0 0 0 C[33]
flabel metal1 30 -2691 438 -2630 1 FreeSans 800 0 0 0 C[34]
flabel metal1 30 -2833 438 -2772 1 FreeSans 800 0 0 0 C[35]
flabel metal1 30 -2975 438 -2914 1 FreeSans 800 0 0 0 C[36]
flabel metal1 30 -3117 438 -3056 1 FreeSans 800 0 0 0 C[37]
flabel metal1 30 -3259 438 -3198 1 FreeSans 800 0 0 0 C[38]
flabel metal1 30 -3401 438 -3340 1 FreeSans 800 0 0 0 C[39]
flabel metal1 30 -3543 438 -3482 1 FreeSans 800 0 0 0 C[40]
flabel metal1 30 -3685 438 -3624 1 FreeSans 800 0 0 0 C[41]
flabel metal1 30 -3827 438 -3766 1 FreeSans 800 0 0 0 C[42]
flabel metal1 30 -3969 438 -3908 1 FreeSans 800 0 0 0 C[43]
flabel metal1 30 -4111 438 -4050 1 FreeSans 800 0 0 0 C[44]
flabel metal1 30 -4253 438 -4192 1 FreeSans 800 0 0 0 C[45]
flabel metal1 30 -4395 438 -4334 1 FreeSans 800 0 0 0 C[46]
flabel metal1 30 -4537 438 -4476 1 FreeSans 800 0 0 0 C[47]
flabel metal1 60835 -138 61307 -77 1 FreeSans 800 0 0 0 C[112]
flabel metal1 60835 -280 61307 -219 1 FreeSans 800 0 0 0 C[113]
flabel metal1 60835 -422 61307 -361 1 FreeSans 800 0 0 0 C[114]
flabel metal1 60835 -564 61307 -503 1 FreeSans 800 0 0 0 C[115]
flabel metal1 60835 -706 61307 -645 1 FreeSans 800 0 0 0 C[116]
flabel metal1 60835 -848 61307 -787 1 FreeSans 800 0 0 0 C[117]
flabel metal1 60835 -990 61307 -929 1 FreeSans 800 0 0 0 C[118]
flabel metal1 60835 -1132 61307 -1071 1 FreeSans 800 0 0 0 C[119]
flabel metal1 60835 -1274 61307 -1213 1 FreeSans 800 0 0 0 C[120]
flabel metal1 60835 -1416 61307 -1355 1 FreeSans 800 0 0 0 C[121]
flabel metal1 60835 -1558 61307 -1497 1 FreeSans 800 0 0 0 C[122]
flabel metal1 60835 -1700 61307 -1639 1 FreeSans 800 0 0 0 C[123]
flabel metal1 60835 -1842 61307 -1781 1 FreeSans 800 0 0 0 C[124]
flabel metal1 60835 -1984 61307 -1923 1 FreeSans 800 0 0 0 C[125]
flabel metal1 60835 -2126 61307 -2065 1 FreeSans 800 0 0 0 C[126]
flabel metal1 60835 -2268 61307 -2207 1 FreeSans 800 0 0 0 C[127]
flabel metal1 60835 -2410 61307 -2349 1 FreeSans 800 0 0 0 C[63]
flabel metal1 60835 -2552 61307 -2491 1 FreeSans 800 0 0 0 C[62]
flabel metal1 60835 -2694 61307 -2633 1 FreeSans 800 0 0 0 C[61]
flabel metal1 60835 -2836 61307 -2775 1 FreeSans 800 0 0 0 C[60]
flabel metal1 60835 -2978 61307 -2917 1 FreeSans 800 0 0 0 C[59]
flabel metal1 60835 -3120 61307 -3059 1 FreeSans 800 0 0 0 C[58]
flabel metal1 60835 -3262 61307 -3201 1 FreeSans 800 0 0 0 C[57]
flabel metal1 60835 -3404 61307 -3343 1 FreeSans 800 0 0 0 C[56]
flabel metal1 60835 -3546 61307 -3485 1 FreeSans 800 0 0 0 C[55]
flabel metal1 60835 -3688 61307 -3627 1 FreeSans 800 0 0 0 C[54]
flabel metal1 60835 -3830 61307 -3769 1 FreeSans 800 0 0 0 C[53]
flabel metal1 60835 -3972 61307 -3911 1 FreeSans 800 0 0 0 C[52]
flabel metal1 60835 -4114 61307 -4053 1 FreeSans 800 0 0 0 C[51]
flabel metal1 60835 -4256 61307 -4195 1 FreeSans 800 0 0 0 C[50]
flabel metal1 60835 -4398 61307 -4337 1 FreeSans 800 0 0 0 C[49]
flabel metal1 60835 -4540 61307 -4479 1 FreeSans 800 0 0 0 C[48]
flabel metal3 -280 -2728 -34 -2638 1 FreeSans 400 0 0 0 RESET
<< end >>
