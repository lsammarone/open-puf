magic
tech sky130A
magscale 1 2
timestamp 1654402208
<< error_p >>
rect 19 181 77 187
rect 19 147 31 181
rect 19 141 77 147
rect -77 -147 -19 -141
rect -77 -181 -65 -147
rect -77 -187 -19 -181
<< nwell >>
rect -65 162 161 200
rect -161 -162 161 162
rect -161 -200 65 -162
<< pmoshvt >>
rect -63 -100 -33 100
rect 33 -100 63 100
<< pdiff >>
rect -125 85 -63 100
rect -125 51 -113 85
rect -79 51 -63 85
rect -125 17 -63 51
rect -125 -17 -113 17
rect -79 -17 -63 17
rect -125 -51 -63 -17
rect -125 -85 -113 -51
rect -79 -85 -63 -51
rect -125 -100 -63 -85
rect -33 85 33 100
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -100 33 -85
rect 63 85 125 100
rect 63 51 79 85
rect 113 51 125 85
rect 63 17 125 51
rect 63 -17 79 17
rect 113 -17 125 17
rect 63 -51 125 -17
rect 63 -85 79 -51
rect 113 -85 125 -51
rect 63 -100 125 -85
<< pdiffc >>
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
<< poly >>
rect 15 181 81 197
rect 15 147 31 181
rect 65 147 81 181
rect 15 131 81 147
rect -63 100 -33 126
rect 33 100 63 131
rect -63 -131 -33 -100
rect 33 -126 63 -100
rect -81 -147 -15 -131
rect -81 -181 -65 -147
rect -31 -181 -15 -147
rect -81 -197 -15 -181
<< polycont >>
rect 31 147 65 181
rect -65 -181 -31 -147
<< locali >>
rect 15 147 31 181
rect 65 147 81 181
rect -113 85 -79 104
rect -113 17 -79 19
rect -113 -19 -79 -17
rect -113 -104 -79 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 79 85 113 104
rect 79 17 113 19
rect 79 -19 113 -17
rect 79 -104 113 -85
rect -81 -181 -65 -147
rect -31 -181 -15 -147
<< viali >>
rect 31 147 65 181
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect -65 -181 -31 -147
<< metal1 >>
rect 19 181 77 187
rect 19 147 31 181
rect 65 147 77 181
rect 19 141 77 147
rect -119 53 -73 100
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -100 -73 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 73 53 119 100
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -100 119 -53
rect -77 -147 -19 -141
rect -77 -181 -65 -147
rect -31 -181 -19 -147
rect -77 -187 -19 -181
<< end >>
