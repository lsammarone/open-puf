magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< locali >>
rect 159 1160 171 1194
rect 205 1160 243 1194
rect 277 1160 315 1194
rect 349 1160 387 1194
rect 421 1160 459 1194
rect 493 1160 505 1194
rect 48 1020 82 1058
rect 48 948 82 986
rect 48 876 82 914
rect 48 804 82 842
rect 48 732 82 770
rect 48 660 82 698
rect 48 588 82 626
rect 48 516 82 554
rect 48 444 82 482
rect 48 372 82 410
rect 48 300 82 338
rect 48 228 82 266
rect 48 122 82 194
rect 582 1020 616 1058
rect 582 948 616 986
rect 582 876 616 914
rect 582 804 616 842
rect 582 732 616 770
rect 582 660 616 698
rect 582 588 616 626
rect 582 516 616 554
rect 582 444 616 482
rect 582 372 616 410
rect 582 300 616 338
rect 582 228 616 266
rect 582 122 616 194
rect 159 20 171 54
rect 205 20 243 54
rect 277 20 315 54
rect 349 20 387 54
rect 421 20 459 54
rect 493 20 505 54
<< viali >>
rect 171 1160 205 1194
rect 243 1160 277 1194
rect 315 1160 349 1194
rect 387 1160 421 1194
rect 459 1160 493 1194
rect 48 1058 82 1092
rect 48 986 82 1020
rect 48 914 82 948
rect 48 842 82 876
rect 48 770 82 804
rect 48 698 82 732
rect 48 626 82 660
rect 48 554 82 588
rect 48 482 82 516
rect 48 410 82 444
rect 48 338 82 372
rect 48 266 82 300
rect 48 194 82 228
rect 582 1058 616 1092
rect 582 986 616 1020
rect 582 914 616 948
rect 582 842 616 876
rect 582 770 616 804
rect 582 698 616 732
rect 582 626 616 660
rect 582 554 616 588
rect 582 482 616 516
rect 582 410 616 444
rect 582 338 616 372
rect 582 266 616 300
rect 582 194 616 228
rect 171 20 205 54
rect 243 20 277 54
rect 315 20 349 54
rect 387 20 421 54
rect 459 20 493 54
<< obsli1 >>
rect 159 98 193 1116
rect 315 98 349 1116
rect 471 98 505 1116
<< metal1 >>
rect 159 1194 505 1214
rect 159 1160 171 1194
rect 205 1160 243 1194
rect 277 1160 315 1194
rect 349 1160 387 1194
rect 421 1160 459 1194
rect 493 1160 505 1194
rect 159 1148 505 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 110 94 194
rect 570 1092 628 1104
rect 570 1058 582 1092
rect 616 1058 628 1092
rect 570 1020 628 1058
rect 570 986 582 1020
rect 616 986 628 1020
rect 570 948 628 986
rect 570 914 582 948
rect 616 914 628 948
rect 570 876 628 914
rect 570 842 582 876
rect 616 842 628 876
rect 570 804 628 842
rect 570 770 582 804
rect 616 770 628 804
rect 570 732 628 770
rect 570 698 582 732
rect 616 698 628 732
rect 570 660 628 698
rect 570 626 582 660
rect 616 626 628 660
rect 570 588 628 626
rect 570 554 582 588
rect 616 554 628 588
rect 570 516 628 554
rect 570 482 582 516
rect 616 482 628 516
rect 570 444 628 482
rect 570 410 582 444
rect 616 410 628 444
rect 570 372 628 410
rect 570 338 582 372
rect 616 338 628 372
rect 570 300 628 338
rect 570 266 582 300
rect 616 266 628 300
rect 570 228 628 266
rect 570 194 582 228
rect 616 194 628 228
rect 570 110 628 194
rect 159 54 505 66
rect 159 20 171 54
rect 205 20 243 54
rect 277 20 315 54
rect 349 20 387 54
rect 421 20 459 54
rect 493 20 505 54
rect 159 0 505 20
<< obsm1 >>
rect 150 110 202 1104
rect 306 110 358 1104
rect 462 110 514 1104
<< metal2 >>
rect 10 632 654 1104
rect 10 110 654 582
<< labels >>
rlabel viali s 582 1058 616 1092 6 BULK
port 1 nsew
rlabel viali s 582 986 616 1020 6 BULK
port 1 nsew
rlabel viali s 582 914 616 948 6 BULK
port 1 nsew
rlabel viali s 582 842 616 876 6 BULK
port 1 nsew
rlabel viali s 582 770 616 804 6 BULK
port 1 nsew
rlabel viali s 582 698 616 732 6 BULK
port 1 nsew
rlabel viali s 582 626 616 660 6 BULK
port 1 nsew
rlabel viali s 582 554 616 588 6 BULK
port 1 nsew
rlabel viali s 582 482 616 516 6 BULK
port 1 nsew
rlabel viali s 582 410 616 444 6 BULK
port 1 nsew
rlabel viali s 582 338 616 372 6 BULK
port 1 nsew
rlabel viali s 582 266 616 300 6 BULK
port 1 nsew
rlabel viali s 582 194 616 228 6 BULK
port 1 nsew
rlabel viali s 48 1058 82 1092 6 BULK
port 1 nsew
rlabel viali s 48 986 82 1020 6 BULK
port 1 nsew
rlabel viali s 48 914 82 948 6 BULK
port 1 nsew
rlabel viali s 48 842 82 876 6 BULK
port 1 nsew
rlabel viali s 48 770 82 804 6 BULK
port 1 nsew
rlabel viali s 48 698 82 732 6 BULK
port 1 nsew
rlabel viali s 48 626 82 660 6 BULK
port 1 nsew
rlabel viali s 48 554 82 588 6 BULK
port 1 nsew
rlabel viali s 48 482 82 516 6 BULK
port 1 nsew
rlabel viali s 48 410 82 444 6 BULK
port 1 nsew
rlabel viali s 48 338 82 372 6 BULK
port 1 nsew
rlabel viali s 48 266 82 300 6 BULK
port 1 nsew
rlabel viali s 48 194 82 228 6 BULK
port 1 nsew
rlabel locali s 582 122 616 1092 6 BULK
port 1 nsew
rlabel locali s 48 122 82 1092 6 BULK
port 1 nsew
rlabel metal1 s 570 110 628 1104 6 BULK
port 1 nsew
rlabel metal1 s 36 110 94 1104 6 BULK
port 1 nsew
rlabel metal2 s 10 632 654 1104 6 DRAIN
port 2 nsew
rlabel viali s 459 1160 493 1194 6 GATE
port 3 nsew
rlabel viali s 459 20 493 54 6 GATE
port 3 nsew
rlabel viali s 387 1160 421 1194 6 GATE
port 3 nsew
rlabel viali s 387 20 421 54 6 GATE
port 3 nsew
rlabel viali s 315 1160 349 1194 6 GATE
port 3 nsew
rlabel viali s 315 20 349 54 6 GATE
port 3 nsew
rlabel viali s 243 1160 277 1194 6 GATE
port 3 nsew
rlabel viali s 243 20 277 54 6 GATE
port 3 nsew
rlabel viali s 171 1160 205 1194 6 GATE
port 3 nsew
rlabel viali s 171 20 205 54 6 GATE
port 3 nsew
rlabel locali s 159 1160 505 1194 6 GATE
port 3 nsew
rlabel locali s 159 20 505 54 6 GATE
port 3 nsew
rlabel metal1 s 159 1148 505 1214 6 GATE
port 3 nsew
rlabel metal1 s 159 0 505 66 6 GATE
port 3 nsew
rlabel metal2 s 10 110 654 582 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 664 1214
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9867544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9851508
<< end >>
