magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 1 21 459 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 343 47 373 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 343 297 373 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 47 163 177
rect 193 47 247 177
rect 277 47 343 177
rect 373 161 433 177
rect 373 127 383 161
rect 417 127 433 161
rect 373 93 433 127
rect 373 59 383 93
rect 417 59 433 93
rect 373 47 433 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 297 247 383
rect 277 485 343 497
rect 277 451 293 485
rect 327 451 343 485
rect 277 417 343 451
rect 277 383 293 417
rect 327 383 343 417
rect 277 349 343 383
rect 277 315 293 349
rect 327 315 343 349
rect 277 297 343 315
rect 373 485 433 497
rect 373 451 383 485
rect 417 451 433 485
rect 373 417 433 451
rect 373 383 383 417
rect 417 383 433 417
rect 373 297 433 383
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 383 127 417 161
rect 383 59 417 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 203 383 237 417
rect 293 451 327 485
rect 293 383 327 417
rect 293 315 327 349
rect 383 451 417 485
rect 383 383 417 417
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 343 497 373 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 343 265 373 297
rect 25 249 109 265
rect 25 215 35 249
rect 69 215 109 249
rect 25 199 109 215
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 151 199 205 215
rect 247 249 301 265
rect 247 215 257 249
rect 291 215 301 249
rect 247 199 301 215
rect 343 249 439 265
rect 343 215 395 249
rect 429 215 439 249
rect 343 199 439 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 343 177 373 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 343 21 373 47
<< polycont >>
rect 35 215 69 249
rect 161 215 195 249
rect 257 215 291 249
rect 395 215 429 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 17 485 69 527
rect 17 451 35 485
rect 17 417 69 451
rect 17 383 35 417
rect 17 349 69 383
rect 17 315 35 349
rect 17 299 69 315
rect 103 485 169 493
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 203 485 237 527
rect 203 417 237 451
rect 203 367 237 383
rect 277 485 343 493
rect 277 451 293 485
rect 327 451 343 485
rect 277 417 343 451
rect 277 383 293 417
rect 327 383 343 417
rect 103 315 119 349
rect 153 333 169 349
rect 277 349 343 383
rect 383 485 439 527
rect 417 451 439 485
rect 383 417 439 451
rect 417 383 439 417
rect 383 367 439 383
rect 277 333 293 349
rect 153 315 293 333
rect 327 333 343 349
rect 327 315 359 333
rect 103 299 359 315
rect 22 249 79 265
rect 22 215 35 249
rect 69 215 79 249
rect 22 199 79 215
rect 119 249 195 265
rect 119 215 161 249
rect 119 199 195 215
rect 229 249 291 265
rect 229 215 257 249
rect 229 199 291 215
rect 18 161 85 165
rect 18 127 35 161
rect 69 127 85 161
rect 18 93 85 127
rect 18 59 35 93
rect 69 59 85 93
rect 119 60 162 199
rect 229 165 270 199
rect 325 165 359 299
rect 395 249 443 333
rect 429 215 443 249
rect 395 199 443 215
rect 200 60 270 165
rect 304 161 443 165
rect 304 127 383 161
rect 417 127 443 161
rect 304 93 443 127
rect 18 17 85 59
rect 304 59 383 93
rect 417 59 443 93
rect 304 51 443 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
flabel locali s 122 221 156 255 0 FreeSans 250 0 0 0 C
port 3 nsew signal input
flabel locali s 214 85 248 119 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 306 85 340 119 0 FreeSans 250 0 0 0 Y
port 9 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 250 0 0 0 D
port 4 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 nand4_1
rlabel metal1 s 0 -48 460 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 460 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 460 544
string GDS_END 1882228
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1877024
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 11.500 0.000 
<< end >>
