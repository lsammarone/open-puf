magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 1 21 1563 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1107 47 1137 177
rect 1191 47 1221 177
rect 1275 47 1305 177
rect 1359 47 1389 177
rect 1443 47 1473 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 755 297 785 497
rect 839 297 869 497
rect 923 297 953 497
rect 1007 297 1037 497
rect 1191 297 1221 497
rect 1275 297 1305 497
rect 1359 297 1389 497
rect 1443 297 1473 497
<< ndiff >>
rect 27 101 79 177
rect 27 67 35 101
rect 69 67 79 101
rect 27 47 79 67
rect 109 93 163 177
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 101 247 177
rect 193 67 203 101
rect 237 67 247 101
rect 193 47 247 67
rect 277 93 331 177
rect 277 59 287 93
rect 321 59 331 93
rect 277 47 331 59
rect 361 101 415 177
rect 361 67 371 101
rect 405 67 415 101
rect 361 47 415 67
rect 445 93 499 177
rect 445 59 455 93
rect 489 59 499 93
rect 445 47 499 59
rect 529 161 583 177
rect 529 127 539 161
rect 573 127 583 161
rect 529 47 583 127
rect 613 93 667 177
rect 613 59 623 93
rect 657 59 667 93
rect 613 47 667 59
rect 697 161 749 177
rect 697 127 707 161
rect 741 127 749 161
rect 697 47 749 127
rect 803 161 855 177
rect 803 127 811 161
rect 845 127 855 161
rect 803 47 855 127
rect 885 93 939 177
rect 885 59 895 93
rect 929 59 939 93
rect 885 47 939 59
rect 969 161 1023 177
rect 969 127 979 161
rect 1013 127 1023 161
rect 969 47 1023 127
rect 1053 93 1107 177
rect 1053 59 1063 93
rect 1097 59 1107 93
rect 1053 47 1107 59
rect 1137 161 1191 177
rect 1137 127 1147 161
rect 1181 127 1191 161
rect 1137 47 1191 127
rect 1221 93 1275 177
rect 1221 59 1231 93
rect 1265 59 1275 93
rect 1221 47 1275 59
rect 1305 101 1359 177
rect 1305 67 1315 101
rect 1349 67 1359 101
rect 1305 47 1359 67
rect 1389 93 1443 177
rect 1389 59 1399 93
rect 1433 59 1443 93
rect 1389 47 1443 59
rect 1473 101 1537 177
rect 1473 67 1483 101
rect 1517 67 1537 101
rect 1473 47 1537 67
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 297 79 375
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 297 163 383
rect 193 477 247 497
rect 193 443 203 477
rect 237 443 247 477
rect 193 409 247 443
rect 193 375 203 409
rect 237 375 247 409
rect 193 297 247 375
rect 277 485 331 497
rect 277 451 287 485
rect 321 451 331 485
rect 277 417 331 451
rect 277 383 287 417
rect 321 383 331 417
rect 277 297 331 383
rect 361 477 415 497
rect 361 443 371 477
rect 405 443 415 477
rect 361 409 415 443
rect 361 375 371 409
rect 405 375 415 409
rect 361 297 415 375
rect 445 485 499 497
rect 445 451 455 485
rect 489 451 499 485
rect 445 417 499 451
rect 445 383 455 417
rect 489 383 499 417
rect 445 297 499 383
rect 529 477 583 497
rect 529 443 539 477
rect 573 443 583 477
rect 529 409 583 443
rect 529 375 539 409
rect 573 375 583 409
rect 529 297 583 375
rect 613 485 667 497
rect 613 451 623 485
rect 657 451 667 485
rect 613 417 667 451
rect 613 383 623 417
rect 657 383 667 417
rect 613 297 667 383
rect 697 477 755 497
rect 697 443 707 477
rect 741 443 755 477
rect 697 409 755 443
rect 697 375 707 409
rect 741 375 755 409
rect 697 297 755 375
rect 785 485 839 497
rect 785 451 795 485
rect 829 451 839 485
rect 785 417 839 451
rect 785 383 795 417
rect 829 383 839 417
rect 785 297 839 383
rect 869 477 923 497
rect 869 443 879 477
rect 913 443 923 477
rect 869 409 923 443
rect 869 375 879 409
rect 913 375 923 409
rect 869 297 923 375
rect 953 485 1007 497
rect 953 451 963 485
rect 997 451 1007 485
rect 953 297 1007 451
rect 1037 477 1191 497
rect 1037 443 1047 477
rect 1081 443 1191 477
rect 1037 377 1191 443
rect 1037 343 1047 377
rect 1081 343 1191 377
rect 1037 297 1191 343
rect 1221 417 1275 497
rect 1221 383 1231 417
rect 1265 383 1275 417
rect 1221 297 1275 383
rect 1305 485 1359 497
rect 1305 451 1315 485
rect 1349 451 1359 485
rect 1305 297 1359 451
rect 1389 417 1443 497
rect 1389 383 1399 417
rect 1433 383 1443 417
rect 1389 297 1443 383
rect 1473 485 1537 497
rect 1473 451 1483 485
rect 1517 451 1537 485
rect 1473 417 1537 451
rect 1473 383 1483 417
rect 1517 383 1537 417
rect 1473 349 1537 383
rect 1473 315 1483 349
rect 1517 315 1537 349
rect 1473 297 1537 315
<< ndiffc >>
rect 35 67 69 101
rect 119 59 153 93
rect 203 67 237 101
rect 287 59 321 93
rect 371 67 405 101
rect 455 59 489 93
rect 539 127 573 161
rect 623 59 657 93
rect 707 127 741 161
rect 811 127 845 161
rect 895 59 929 93
rect 979 127 1013 161
rect 1063 59 1097 93
rect 1147 127 1181 161
rect 1231 59 1265 93
rect 1315 67 1349 101
rect 1399 59 1433 93
rect 1483 67 1517 101
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 451 153 485
rect 119 383 153 417
rect 203 443 237 477
rect 203 375 237 409
rect 287 451 321 485
rect 287 383 321 417
rect 371 443 405 477
rect 371 375 405 409
rect 455 451 489 485
rect 455 383 489 417
rect 539 443 573 477
rect 539 375 573 409
rect 623 451 657 485
rect 623 383 657 417
rect 707 443 741 477
rect 707 375 741 409
rect 795 451 829 485
rect 795 383 829 417
rect 879 443 913 477
rect 879 375 913 409
rect 963 451 997 485
rect 1047 443 1081 477
rect 1047 343 1081 377
rect 1231 383 1265 417
rect 1315 451 1349 485
rect 1399 383 1433 417
rect 1483 451 1517 485
rect 1483 383 1517 417
rect 1483 315 1517 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 755 497 785 523
rect 839 497 869 523
rect 923 497 953 523
rect 1007 497 1037 523
rect 1191 497 1221 523
rect 1275 497 1305 523
rect 1359 497 1389 523
rect 1443 497 1473 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 22 249 361 265
rect 22 215 40 249
rect 74 215 114 249
rect 148 215 188 249
rect 222 215 262 249
rect 296 215 361 249
rect 22 199 361 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 415 265 445 297
rect 499 265 529 297
rect 583 265 613 297
rect 667 265 697 297
rect 415 249 697 265
rect 415 215 425 249
rect 459 215 499 249
rect 533 215 573 249
rect 607 215 647 249
rect 681 215 697 249
rect 415 199 697 215
rect 755 269 785 297
rect 839 269 869 297
rect 923 269 953 297
rect 1007 269 1037 297
rect 755 265 1037 269
rect 1191 265 1221 297
rect 1275 265 1305 297
rect 1359 265 1389 297
rect 1443 265 1473 297
rect 755 249 1137 265
rect 755 215 765 249
rect 799 215 839 249
rect 873 215 913 249
rect 947 215 987 249
rect 1021 215 1137 249
rect 755 202 1137 215
rect 755 199 1053 202
rect 415 177 445 199
rect 499 177 529 199
rect 583 177 613 199
rect 667 177 697 199
rect 855 177 885 199
rect 939 177 969 199
rect 1023 177 1053 199
rect 1107 177 1137 202
rect 1179 249 1473 265
rect 1179 215 1189 249
rect 1223 215 1263 249
rect 1297 215 1337 249
rect 1371 215 1473 249
rect 1179 199 1473 215
rect 1191 177 1221 199
rect 1275 177 1305 199
rect 1359 177 1389 199
rect 1443 177 1473 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1107 21 1137 47
rect 1191 21 1221 47
rect 1275 21 1305 47
rect 1359 21 1389 47
rect 1443 21 1473 47
<< polycont >>
rect 40 215 74 249
rect 114 215 148 249
rect 188 215 222 249
rect 262 215 296 249
rect 425 215 459 249
rect 499 215 533 249
rect 573 215 607 249
rect 647 215 681 249
rect 765 215 799 249
rect 839 215 873 249
rect 913 215 947 249
rect 987 215 1021 249
rect 1189 215 1223 249
rect 1263 215 1297 249
rect 1337 215 1371 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 35 477 69 493
rect 35 409 69 443
rect 103 485 169 527
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 203 477 237 493
rect 203 409 237 443
rect 35 333 69 375
rect 271 485 337 527
rect 271 451 287 485
rect 321 451 337 485
rect 271 417 337 451
rect 271 383 287 417
rect 321 383 337 417
rect 371 477 405 493
rect 371 409 405 443
rect 203 333 237 375
rect 439 485 505 527
rect 439 451 455 485
rect 489 451 505 485
rect 439 417 505 451
rect 439 383 455 417
rect 489 383 505 417
rect 539 477 573 493
rect 539 409 573 443
rect 371 333 405 375
rect 607 485 673 527
rect 607 451 623 485
rect 657 451 673 485
rect 607 417 673 451
rect 607 383 623 417
rect 657 383 673 417
rect 707 477 741 493
rect 707 409 741 443
rect 539 333 573 375
rect 779 485 845 527
rect 779 451 795 485
rect 829 451 845 485
rect 779 417 845 451
rect 779 383 795 417
rect 829 383 845 417
rect 879 477 913 493
rect 947 485 1013 527
rect 947 451 963 485
rect 997 451 1013 485
rect 1047 485 1081 493
rect 1047 477 1315 485
rect 879 409 913 443
rect 707 333 741 375
rect 879 333 913 375
rect 1081 451 1315 477
rect 1349 451 1483 485
rect 1517 451 1533 485
rect 1047 377 1081 443
rect 1483 417 1533 451
rect 1215 383 1231 417
rect 1265 383 1399 417
rect 1433 383 1449 417
rect 1047 333 1081 343
rect 35 299 1081 333
rect 24 249 347 265
rect 24 215 40 249
rect 74 215 114 249
rect 148 215 188 249
rect 222 215 262 249
rect 296 215 347 249
rect 24 199 347 215
rect 387 249 710 265
rect 387 215 425 249
rect 459 215 499 249
rect 533 215 573 249
rect 607 215 647 249
rect 681 215 710 249
rect 387 199 710 215
rect 765 249 1084 265
rect 799 215 839 249
rect 873 215 913 249
rect 947 215 987 249
rect 1021 215 1084 249
rect 765 199 1084 215
rect 1134 249 1371 326
rect 1134 215 1189 249
rect 1223 215 1263 249
rect 1297 215 1337 249
rect 1134 199 1371 215
rect 1409 161 1449 383
rect 1517 383 1533 417
rect 1483 349 1533 383
rect 1517 315 1533 349
rect 1483 299 1533 315
rect 35 127 539 161
rect 573 127 707 161
rect 741 127 757 161
rect 795 127 811 161
rect 845 127 979 161
rect 1013 127 1147 161
rect 1181 127 1517 161
rect 35 101 69 127
rect 203 101 237 127
rect 35 51 69 67
rect 103 59 119 93
rect 153 59 169 93
rect 103 17 169 59
rect 371 101 405 127
rect 203 51 237 67
rect 271 59 287 93
rect 321 59 337 93
rect 271 17 337 59
rect 1315 101 1349 127
rect 371 51 405 67
rect 439 59 455 93
rect 489 59 623 93
rect 657 59 895 93
rect 929 59 1063 93
rect 1097 59 1113 93
rect 1215 59 1231 93
rect 1265 59 1281 93
rect 1215 17 1281 59
rect 1483 101 1517 127
rect 1315 51 1349 67
rect 1383 59 1399 93
rect 1433 59 1449 93
rect 1383 17 1449 59
rect 1483 51 1517 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel locali s 1414 153 1448 187 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1414 221 1448 255 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1414 289 1448 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1414 357 1448 391 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1138 289 1172 323 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 770 221 804 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1138 221 1172 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1322 289 1356 323 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1230 289 1264 323 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1322 221 1356 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1230 221 1264 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 1046 221 1080 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 674 221 708 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 954 221 988 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 862 221 896 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 a31oi_4
rlabel metal1 s 0 -48 1564 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1564 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_END 4164820
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4151954
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 39.100 0.000 
<< end >>
