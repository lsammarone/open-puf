magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 21 905 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 363 47 393 177
rect 466 47 496 177
rect 567 47 597 177
rect 667 47 697 177
rect 767 47 797 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 315 297 345 497
rect 466 297 496 497
rect 567 297 597 497
rect 667 297 697 497
rect 767 297 797 497
<< ndiff >>
rect 27 161 79 177
rect 27 127 35 161
rect 69 127 79 161
rect 27 93 79 127
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 161 163 177
rect 109 127 119 161
rect 153 127 163 161
rect 109 93 163 127
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 161 245 177
rect 193 127 203 161
rect 237 127 245 161
rect 193 93 245 127
rect 193 59 203 93
rect 237 59 245 93
rect 193 47 245 59
rect 299 161 363 177
rect 299 127 307 161
rect 341 127 363 161
rect 299 93 363 127
rect 299 59 307 93
rect 341 59 363 93
rect 299 47 363 59
rect 393 161 466 177
rect 393 127 413 161
rect 447 127 466 161
rect 393 93 466 127
rect 393 59 413 93
rect 447 59 466 93
rect 393 47 466 59
rect 496 93 567 177
rect 496 59 506 93
rect 540 59 567 93
rect 496 47 567 59
rect 597 161 667 177
rect 597 127 607 161
rect 641 127 667 161
rect 597 93 667 127
rect 597 59 607 93
rect 641 59 667 93
rect 597 47 667 59
rect 697 93 767 177
rect 697 59 711 93
rect 745 59 767 93
rect 697 47 767 59
rect 797 161 879 177
rect 797 127 829 161
rect 863 127 879 161
rect 797 93 879 127
rect 797 59 829 93
rect 863 59 879 93
rect 797 47 879 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 315 497
rect 193 383 203 485
rect 305 383 315 485
rect 193 349 315 383
rect 193 315 203 349
rect 237 315 315 349
rect 193 297 315 315
rect 345 485 466 497
rect 345 451 355 485
rect 389 451 466 485
rect 345 417 466 451
rect 345 383 355 417
rect 389 383 466 417
rect 345 349 466 383
rect 345 315 355 349
rect 389 315 466 349
rect 345 297 466 315
rect 496 297 567 497
rect 597 297 667 497
rect 697 297 767 497
rect 797 485 879 497
rect 797 451 829 485
rect 863 451 879 485
rect 797 417 879 451
rect 797 383 829 417
rect 863 383 879 417
rect 797 349 879 383
rect 797 315 829 349
rect 863 315 879 349
rect 797 297 879 315
<< ndiffc >>
rect 35 127 69 161
rect 35 59 69 93
rect 119 127 153 161
rect 119 59 153 93
rect 203 127 237 161
rect 203 59 237 93
rect 307 127 341 161
rect 307 59 341 93
rect 413 127 447 161
rect 413 59 447 93
rect 506 59 540 93
rect 607 127 641 161
rect 607 59 641 93
rect 711 59 745 93
rect 829 127 863 161
rect 829 59 863 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 383 305 485
rect 203 315 237 349
rect 355 451 389 485
rect 355 383 389 417
rect 355 315 389 349
rect 829 451 863 485
rect 829 383 863 417
rect 829 315 863 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 315 497 345 523
rect 466 497 496 523
rect 567 497 597 523
rect 667 497 697 523
rect 767 497 797 523
rect 79 269 109 297
rect 163 269 193 297
rect 79 259 193 269
rect 315 259 345 297
rect 466 265 496 297
rect 567 265 597 297
rect 667 265 697 297
rect 767 265 797 297
rect 79 249 259 259
rect 79 215 209 249
rect 243 215 259 249
rect 79 205 259 215
rect 315 249 421 259
rect 315 215 371 249
rect 405 215 421 249
rect 315 205 421 215
rect 466 249 525 265
rect 466 215 481 249
rect 515 215 525 249
rect 79 195 193 205
rect 79 177 109 195
rect 163 177 193 195
rect 363 177 393 205
rect 466 199 525 215
rect 567 249 625 265
rect 567 215 581 249
rect 615 215 625 249
rect 567 199 625 215
rect 667 249 725 265
rect 667 215 681 249
rect 715 215 725 249
rect 667 199 725 215
rect 767 249 825 265
rect 767 215 781 249
rect 815 215 825 249
rect 767 199 825 215
rect 466 177 496 199
rect 567 177 597 199
rect 667 177 697 199
rect 767 177 797 199
rect 79 21 109 47
rect 163 21 193 47
rect 363 21 393 47
rect 466 21 496 47
rect 567 21 597 47
rect 667 21 697 47
rect 767 21 797 47
<< polycont >>
rect 209 215 243 249
rect 371 215 405 249
rect 481 215 515 249
rect 581 215 615 249
rect 681 215 715 249
rect 781 215 815 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 17 485 69 527
rect 17 451 35 485
rect 17 417 69 451
rect 17 383 35 417
rect 17 349 69 383
rect 17 315 35 349
rect 17 299 69 315
rect 103 485 169 493
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 103 315 119 349
rect 153 315 169 349
rect 103 299 169 315
rect 203 485 305 527
rect 203 367 305 383
rect 339 485 429 493
rect 339 451 355 485
rect 389 451 429 485
rect 813 485 879 527
rect 339 417 429 451
rect 339 383 355 417
rect 389 383 429 417
rect 203 349 237 367
rect 339 349 429 383
rect 339 333 355 349
rect 203 299 237 315
rect 271 315 355 333
rect 389 315 429 349
rect 271 299 429 315
rect 17 161 69 177
rect 17 127 35 161
rect 17 93 69 127
rect 17 59 35 93
rect 17 17 69 59
rect 103 176 158 299
rect 271 265 320 299
rect 192 249 320 265
rect 192 215 209 249
rect 243 215 320 249
rect 355 249 431 265
rect 355 215 371 249
rect 405 215 431 249
rect 465 249 531 468
rect 465 215 481 249
rect 515 215 531 249
rect 565 249 631 468
rect 565 215 581 249
rect 615 215 631 249
rect 665 249 731 467
rect 813 451 829 485
rect 863 451 879 485
rect 813 417 879 451
rect 813 383 829 417
rect 863 383 879 417
rect 813 349 879 383
rect 813 315 829 349
rect 863 315 879 349
rect 813 299 879 315
rect 665 215 681 249
rect 715 215 731 249
rect 765 249 903 265
rect 765 215 781 249
rect 815 215 903 249
rect 103 161 169 176
rect 103 127 119 161
rect 153 127 169 161
rect 103 93 169 127
rect 103 59 119 93
rect 153 59 169 93
rect 103 51 169 59
rect 203 161 252 177
rect 237 127 252 161
rect 203 93 252 127
rect 237 59 252 93
rect 203 17 252 59
rect 286 170 320 215
rect 286 161 357 170
rect 286 127 307 161
rect 341 127 357 161
rect 286 93 357 127
rect 286 59 307 93
rect 341 59 357 93
rect 286 51 357 59
rect 397 161 879 181
rect 397 127 413 161
rect 447 143 607 161
rect 447 127 463 143
rect 397 93 463 127
rect 591 127 607 143
rect 641 143 829 161
rect 641 127 657 143
rect 397 59 413 93
rect 447 59 463 93
rect 397 51 463 59
rect 497 93 550 109
rect 497 59 506 93
rect 540 59 550 93
rect 497 17 550 59
rect 591 93 657 127
rect 813 127 829 143
rect 863 127 879 161
rect 591 59 607 93
rect 641 59 657 93
rect 591 51 657 59
rect 701 93 755 109
rect 701 59 711 93
rect 745 59 755 93
rect 701 17 755 59
rect 813 93 879 127
rect 813 59 829 93
rect 863 59 879 93
rect 813 51 879 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 857 221 891 255 0 FreeSans 250 0 0 0 A1
port 1 nsew signal input
flabel locali s 673 221 707 255 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 673 289 707 323 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 673 357 707 391 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 673 425 707 459 0 FreeSans 250 0 0 0 A2
port 2 nsew signal input
flabel locali s 581 425 615 459 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 581 357 615 391 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 581 289 615 323 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 250 0 0 0 A3
port 3 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 250 0 0 0 A4
port 4 nsew signal input
flabel locali s 489 289 523 323 0 FreeSans 250 0 0 0 A4
port 4 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 250 0 0 0 B1
port 5 nsew signal input
flabel locali s 122 85 156 119 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel locali s 122 153 156 187 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel locali s 122 221 156 255 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel locali s 122 289 156 323 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel locali s 122 357 156 391 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel locali s 122 425 156 459 0 FreeSans 250 0 0 0 X
port 10 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o41a_2
rlabel metal1 s 0 -48 920 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 708084
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 699004
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 4.600 0.000 
<< end >>
