magic
tech sky130A
magscale 1 2
timestamp 1648127584
<< pwell >>
rect 15 163 615 817
<< nmoslvt >>
rect 171 189 201 791
rect 257 189 287 791
rect 343 189 373 791
rect 429 189 459 791
<< ndiff >>
rect 111 779 171 791
rect 111 745 126 779
rect 160 745 171 779
rect 111 711 171 745
rect 111 677 126 711
rect 160 677 171 711
rect 111 643 171 677
rect 111 609 126 643
rect 160 609 171 643
rect 111 575 171 609
rect 111 541 126 575
rect 160 541 171 575
rect 111 507 171 541
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 779 257 791
rect 201 513 212 779
rect 246 513 257 779
rect 201 467 257 513
rect 201 201 212 467
rect 246 201 257 467
rect 201 189 257 201
rect 287 779 343 791
rect 287 513 298 779
rect 332 513 343 779
rect 287 467 343 513
rect 287 201 298 467
rect 332 201 343 467
rect 287 189 343 201
rect 373 779 429 791
rect 373 513 384 779
rect 418 513 429 779
rect 373 467 429 513
rect 373 201 384 467
rect 418 201 429 467
rect 373 189 429 201
rect 459 779 519 791
rect 459 745 470 779
rect 504 745 519 779
rect 459 711 519 745
rect 459 677 470 711
rect 504 677 519 711
rect 459 643 519 677
rect 459 609 470 643
rect 504 609 519 643
rect 459 575 519 609
rect 459 541 470 575
rect 504 541 519 575
rect 459 507 519 541
rect 459 473 470 507
rect 504 473 519 507
rect 459 439 519 473
rect 459 405 470 439
rect 504 405 519 439
rect 459 371 519 405
rect 459 337 470 371
rect 504 337 519 371
rect 459 303 519 337
rect 459 269 470 303
rect 504 269 519 303
rect 459 235 519 269
rect 459 201 470 235
rect 504 201 519 235
rect 459 189 519 201
<< ndiffc >>
rect 126 745 160 779
rect 126 677 160 711
rect 126 609 160 643
rect 126 541 160 575
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 513 246 779
rect 212 201 246 467
rect 298 513 332 779
rect 298 201 332 467
rect 384 513 418 779
rect 384 201 418 467
rect 470 745 504 779
rect 470 677 504 711
rect 470 609 504 643
rect 470 541 504 575
rect 470 473 504 507
rect 470 405 504 439
rect 470 337 504 371
rect 470 269 504 303
rect 470 201 504 235
<< psubdiff >>
rect 41 779 111 791
rect 41 745 58 779
rect 92 745 111 779
rect 41 711 111 745
rect 41 677 58 711
rect 92 677 111 711
rect 41 643 111 677
rect 41 609 58 643
rect 92 609 111 643
rect 41 575 111 609
rect 41 541 58 575
rect 92 541 111 575
rect 41 507 111 541
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 519 779 589 791
rect 519 745 538 779
rect 572 745 589 779
rect 519 711 589 745
rect 519 677 538 711
rect 572 677 589 711
rect 519 643 589 677
rect 519 609 538 643
rect 572 609 589 643
rect 519 575 589 609
rect 519 541 538 575
rect 572 541 589 575
rect 519 507 589 541
rect 519 473 538 507
rect 572 473 589 507
rect 519 439 589 473
rect 519 405 538 439
rect 572 405 589 439
rect 519 371 589 405
rect 519 337 538 371
rect 572 337 589 371
rect 519 303 589 337
rect 519 269 538 303
rect 572 269 589 303
rect 519 235 589 269
rect 519 201 538 235
rect 572 201 589 235
rect 519 189 589 201
<< psubdiffcont >>
rect 58 745 92 779
rect 58 677 92 711
rect 58 609 92 643
rect 58 541 92 575
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 538 745 572 779
rect 538 677 572 711
rect 538 609 572 643
rect 538 541 572 575
rect 538 473 572 507
rect 538 405 572 439
rect 538 337 572 371
rect 538 269 572 303
rect 538 201 572 235
<< poly >>
rect 243 891 387 907
rect 120 867 201 883
rect 120 833 136 867
rect 170 833 201 867
rect 243 857 264 891
rect 366 857 387 891
rect 243 841 387 857
rect 429 867 510 883
rect 120 817 201 833
rect 171 791 201 817
rect 257 791 287 841
rect 343 791 373 841
rect 429 833 460 867
rect 494 833 510 867
rect 429 817 510 833
rect 429 791 459 817
rect 171 163 201 189
rect 120 147 201 163
rect 120 113 136 147
rect 170 113 201 147
rect 257 139 287 189
rect 343 139 373 189
rect 429 163 459 189
rect 429 147 510 163
rect 120 97 201 113
rect 243 123 387 139
rect 243 89 264 123
rect 366 89 387 123
rect 429 113 460 147
rect 494 113 510 147
rect 429 97 510 113
rect 243 73 387 89
<< polycont >>
rect 136 833 170 867
rect 264 857 366 891
rect 460 833 494 867
rect 136 113 170 147
rect 264 89 366 123
rect 460 113 494 147
<< locali >>
rect 248 961 382 980
rect 120 867 186 883
rect 120 833 136 867
rect 170 833 186 867
rect 248 855 262 961
rect 368 855 382 961
rect 248 841 382 855
rect 444 867 510 883
rect 120 817 186 833
rect 444 833 460 867
rect 494 833 510 867
rect 444 817 510 833
rect 120 795 160 817
rect 470 795 510 817
rect 41 779 160 795
rect 41 745 58 779
rect 92 759 126 779
rect 94 745 126 759
rect 41 725 60 745
rect 94 725 160 745
rect 41 711 160 725
rect 41 677 58 711
rect 92 687 126 711
rect 94 677 126 687
rect 41 653 60 677
rect 94 653 160 677
rect 41 643 160 653
rect 41 609 58 643
rect 92 615 126 643
rect 94 609 126 615
rect 41 581 60 609
rect 94 581 160 609
rect 41 575 160 581
rect 41 541 58 575
rect 92 543 126 575
rect 94 541 126 543
rect 41 509 60 541
rect 94 509 160 541
rect 41 507 160 509
rect 41 473 58 507
rect 92 473 126 507
rect 41 471 160 473
rect 41 439 60 471
rect 94 439 160 471
rect 41 405 58 439
rect 94 437 126 439
rect 92 405 126 437
rect 41 399 160 405
rect 41 371 60 399
rect 94 371 160 399
rect 41 337 58 371
rect 94 365 126 371
rect 92 337 126 365
rect 41 327 160 337
rect 41 303 60 327
rect 94 303 160 327
rect 41 269 58 303
rect 94 293 126 303
rect 92 269 126 293
rect 41 255 160 269
rect 41 235 60 255
rect 94 235 160 255
rect 41 201 58 235
rect 94 221 126 235
rect 92 201 126 221
rect 41 185 160 201
rect 212 779 246 795
rect 212 471 246 509
rect 212 185 246 201
rect 298 779 332 795
rect 298 471 332 509
rect 298 185 332 201
rect 384 779 418 795
rect 384 471 418 509
rect 384 185 418 201
rect 470 779 589 795
rect 504 759 538 779
rect 504 745 536 759
rect 572 745 589 779
rect 470 725 536 745
rect 570 725 589 745
rect 470 711 589 725
rect 504 687 538 711
rect 504 677 536 687
rect 572 677 589 711
rect 470 653 536 677
rect 570 653 589 677
rect 470 643 589 653
rect 504 615 538 643
rect 504 609 536 615
rect 572 609 589 643
rect 470 581 536 609
rect 570 581 589 609
rect 470 575 589 581
rect 504 543 538 575
rect 504 541 536 543
rect 572 541 589 575
rect 470 509 536 541
rect 570 509 589 541
rect 470 507 589 509
rect 504 473 538 507
rect 572 473 589 507
rect 470 471 589 473
rect 470 439 536 471
rect 570 439 589 471
rect 504 437 536 439
rect 504 405 538 437
rect 572 405 589 439
rect 470 399 589 405
rect 470 371 536 399
rect 570 371 589 399
rect 504 365 536 371
rect 504 337 538 365
rect 572 337 589 371
rect 470 327 589 337
rect 470 303 536 327
rect 570 303 589 327
rect 504 293 536 303
rect 504 269 538 293
rect 572 269 589 303
rect 470 255 589 269
rect 470 235 536 255
rect 570 235 589 255
rect 504 221 536 235
rect 504 201 538 221
rect 572 201 589 235
rect 470 185 589 201
rect 120 163 160 185
rect 470 163 510 185
rect 120 147 186 163
rect 120 113 136 147
rect 170 113 186 147
rect 444 147 510 163
rect 120 97 186 113
rect 248 125 382 139
rect 248 19 262 125
rect 368 19 382 125
rect 444 113 460 147
rect 494 113 510 147
rect 444 97 510 113
rect 248 0 382 19
<< viali >>
rect 262 891 368 961
rect 262 857 264 891
rect 264 857 366 891
rect 366 857 368 891
rect 262 855 368 857
rect 60 745 92 759
rect 92 745 94 759
rect 60 725 94 745
rect 60 677 92 687
rect 92 677 94 687
rect 60 653 94 677
rect 60 609 92 615
rect 92 609 94 615
rect 60 581 94 609
rect 60 541 92 543
rect 92 541 94 543
rect 60 509 94 541
rect 60 439 94 471
rect 60 437 92 439
rect 92 437 94 439
rect 60 371 94 399
rect 60 365 92 371
rect 92 365 94 371
rect 60 303 94 327
rect 60 293 92 303
rect 92 293 94 303
rect 60 235 94 255
rect 60 221 92 235
rect 92 221 94 235
rect 212 725 246 759
rect 212 653 246 687
rect 212 581 246 615
rect 212 513 246 543
rect 212 509 246 513
rect 212 467 246 471
rect 212 437 246 467
rect 212 365 246 399
rect 212 293 246 327
rect 212 221 246 255
rect 298 725 332 759
rect 298 653 332 687
rect 298 581 332 615
rect 298 513 332 543
rect 298 509 332 513
rect 298 467 332 471
rect 298 437 332 467
rect 298 365 332 399
rect 298 293 332 327
rect 298 221 332 255
rect 384 725 418 759
rect 384 653 418 687
rect 384 581 418 615
rect 384 513 418 543
rect 384 509 418 513
rect 384 467 418 471
rect 384 437 418 467
rect 384 365 418 399
rect 384 293 418 327
rect 384 221 418 255
rect 536 745 538 759
rect 538 745 570 759
rect 536 725 570 745
rect 536 677 538 687
rect 538 677 570 687
rect 536 653 570 677
rect 536 609 538 615
rect 538 609 570 615
rect 536 581 570 609
rect 536 541 538 543
rect 538 541 570 543
rect 536 509 570 541
rect 536 439 570 471
rect 536 437 538 439
rect 538 437 570 439
rect 536 371 570 399
rect 536 365 538 371
rect 538 365 570 371
rect 536 303 570 327
rect 536 293 538 303
rect 538 293 570 303
rect 536 235 570 255
rect 536 221 538 235
rect 538 221 570 235
rect 262 123 368 125
rect 262 89 264 123
rect 264 89 366 123
rect 366 89 368 123
rect 262 19 368 89
<< metal1 >>
rect 250 961 380 980
rect 250 855 262 961
rect 368 855 380 961
rect 250 843 380 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 203 759 255 771
rect 203 725 212 759
rect 246 725 255 759
rect 203 687 255 725
rect 203 653 212 687
rect 246 653 255 687
rect 203 615 255 653
rect 203 581 212 615
rect 246 581 255 615
rect 203 543 255 581
rect 203 509 212 543
rect 246 509 255 543
rect 203 471 255 509
rect 203 459 212 471
rect 246 459 255 471
rect 203 399 255 407
rect 203 395 212 399
rect 246 395 255 399
rect 203 331 255 343
rect 203 267 255 279
rect 203 209 255 215
rect 289 765 341 771
rect 289 701 341 713
rect 289 637 341 649
rect 289 581 298 585
rect 332 581 341 585
rect 289 573 341 581
rect 289 509 298 521
rect 332 509 341 521
rect 289 471 341 509
rect 289 437 298 471
rect 332 437 341 471
rect 289 399 341 437
rect 289 365 298 399
rect 332 365 341 399
rect 289 327 341 365
rect 289 293 298 327
rect 332 293 341 327
rect 289 255 341 293
rect 289 221 298 255
rect 332 221 341 255
rect 289 209 341 221
rect 375 759 427 771
rect 375 725 384 759
rect 418 725 427 759
rect 375 687 427 725
rect 375 653 384 687
rect 418 653 427 687
rect 375 615 427 653
rect 375 581 384 615
rect 418 581 427 615
rect 375 543 427 581
rect 375 509 384 543
rect 418 509 427 543
rect 375 471 427 509
rect 375 459 384 471
rect 418 459 427 471
rect 375 399 427 407
rect 375 395 384 399
rect 418 395 427 399
rect 375 331 427 343
rect 375 267 427 279
rect 375 209 427 215
rect 530 759 589 771
rect 530 725 536 759
rect 570 725 589 759
rect 530 687 589 725
rect 530 653 536 687
rect 570 653 589 687
rect 530 615 589 653
rect 530 581 536 615
rect 570 581 589 615
rect 530 543 589 581
rect 530 509 536 543
rect 570 509 589 543
rect 530 471 589 509
rect 530 437 536 471
rect 570 437 589 471
rect 530 399 589 437
rect 530 365 536 399
rect 570 365 589 399
rect 530 327 589 365
rect 530 293 536 327
rect 570 293 589 327
rect 530 255 589 293
rect 530 221 536 255
rect 570 221 589 255
rect 530 209 589 221
rect 250 125 380 137
rect 250 19 262 125
rect 368 19 380 125
rect 250 0 380 19
<< via1 >>
rect 203 437 212 459
rect 212 437 246 459
rect 246 437 255 459
rect 203 407 255 437
rect 203 365 212 395
rect 212 365 246 395
rect 246 365 255 395
rect 203 343 255 365
rect 203 327 255 331
rect 203 293 212 327
rect 212 293 246 327
rect 246 293 255 327
rect 203 279 255 293
rect 203 255 255 267
rect 203 221 212 255
rect 212 221 246 255
rect 246 221 255 255
rect 203 215 255 221
rect 289 759 341 765
rect 289 725 298 759
rect 298 725 332 759
rect 332 725 341 759
rect 289 713 341 725
rect 289 687 341 701
rect 289 653 298 687
rect 298 653 332 687
rect 332 653 341 687
rect 289 649 341 653
rect 289 615 341 637
rect 289 585 298 615
rect 298 585 332 615
rect 332 585 341 615
rect 289 543 341 573
rect 289 521 298 543
rect 298 521 332 543
rect 332 521 341 543
rect 375 437 384 459
rect 384 437 418 459
rect 418 437 427 459
rect 375 407 427 437
rect 375 365 384 395
rect 384 365 418 395
rect 418 365 427 395
rect 375 343 427 365
rect 375 327 427 331
rect 375 293 384 327
rect 384 293 418 327
rect 418 293 427 327
rect 375 279 427 293
rect 375 255 427 267
rect 375 221 384 255
rect 384 221 418 255
rect 418 221 427 255
rect 375 215 427 221
<< metal2 >>
rect 14 765 616 771
rect 14 713 289 765
rect 341 713 616 765
rect 14 701 616 713
rect 14 649 289 701
rect 341 649 616 701
rect 14 637 616 649
rect 14 585 289 637
rect 341 585 616 637
rect 14 573 616 585
rect 14 521 289 573
rect 341 521 616 573
rect 14 515 616 521
rect 14 459 616 465
rect 14 407 203 459
rect 255 407 375 459
rect 427 407 616 459
rect 14 395 616 407
rect 14 343 203 395
rect 255 343 375 395
rect 427 343 616 395
rect 14 331 616 343
rect 14 279 203 331
rect 255 279 375 331
rect 427 279 616 331
rect 14 267 616 279
rect 14 215 203 267
rect 255 215 375 267
rect 427 215 616 267
rect 14 209 616 215
<< labels >>
flabel comment s 182 525 182 525 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 442 520 442 520 0 FreeSans 180 90 0 0 dummy_poly
flabel metal1 s 255 44 374 95 0 FreeSans 200 0 0 0 GATE
port 1 nsew
flabel metal1 s 255 880 374 931 0 FreeSans 200 0 0 0 GATE
port 1 nsew
flabel metal1 s 41 466 100 496 0 FreeSans 200 90 0 0 SUBSTRATE
port 2 nsew
flabel metal1 s 530 469 589 499 0 FreeSans 200 90 0 0 SUBSTRATE
port 2 nsew
flabel metal2 s 14 280 35 408 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal2 s 14 589 35 717 7 FreeSans 300 180 0 0 DRAIN
port 4 nsew
<< properties >>
string GDS_END 6550204
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6537340
<< end >>
