magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1027 203
rect 30 -17 64 21
<< locali >>
rect 28 215 248 255
<< obsli1 >>
rect 0 527 1104 561
rect 19 323 85 493
rect 119 367 153 527
rect 187 323 253 493
rect 287 367 321 527
rect 371 323 405 493
rect 439 367 505 527
rect 539 323 573 493
rect 607 367 673 527
rect 707 323 741 493
rect 775 367 841 527
rect 875 323 909 493
rect 19 289 319 323
rect 371 289 909 323
rect 943 297 1009 527
rect 284 249 319 289
rect 858 263 909 289
rect 284 215 809 249
rect 284 181 319 215
rect 858 211 974 263
rect 858 181 909 211
rect 35 147 319 181
rect 371 147 909 181
rect 35 51 69 147
rect 103 17 169 113
rect 203 52 237 147
rect 271 17 337 113
rect 371 51 405 147
rect 439 17 505 113
rect 539 51 573 147
rect 607 17 673 113
rect 707 51 741 147
rect 775 17 841 113
rect 875 51 909 147
rect 943 17 1009 177
rect 0 -17 1104 17
<< obsm1 >>
rect 0 570 1104 592
rect 0 518 1168 570
rect 0 496 1104 518
rect 404 252 532 264
rect 849 252 979 261
rect 404 224 979 252
rect 404 212 532 224
rect 849 215 979 224
rect 0 26 1104 48
rect 0 -26 1168 26
rect 0 -48 1104 -26
<< metal2 >>
rect 378 210 387 266
rect 443 210 467 266
rect 523 210 532 266
<< via2 >>
rect 387 210 443 266
rect 467 210 523 266
<< obsm2 >>
rect 1027 516 1181 572
rect 1027 -28 1181 28
<< metal3 >>
rect 1026 576 1182 577
rect 1026 512 1032 576
rect 1096 512 1112 576
rect 1176 512 1182 576
rect 1026 511 1182 512
rect 377 270 533 271
rect 377 206 383 270
rect 447 206 463 270
rect 527 206 533 270
rect 377 205 533 206
rect 1026 32 1182 33
rect 1026 -32 1032 32
rect 1096 -32 1112 32
rect 1176 -32 1182 32
rect 1026 -33 1182 -32
<< obsm3 >>
rect -143 206 13 270
<< via3 >>
rect 1032 512 1096 576
rect 1112 512 1176 576
rect 383 266 447 270
rect 383 210 387 266
rect 387 210 443 266
rect 443 210 447 266
rect 383 206 447 210
rect 463 266 527 270
rect 463 210 467 266
rect 467 210 523 266
rect 523 210 527 266
rect 463 206 527 210
rect 1032 -32 1096 32
rect 1112 -32 1176 32
<< metal4 >>
rect 986 576 1222 723
rect 986 512 1032 576
rect 1096 512 1112 576
rect 1176 512 1222 576
rect 986 487 1222 512
rect 292 270 528 390
rect 292 206 383 270
rect 447 206 463 270
rect 527 206 528 270
rect 292 154 528 206
rect 986 32 1222 57
rect 986 -32 1032 32
rect 1096 -32 1112 32
rect 1176 -32 1222 32
rect 986 -179 1222 -32
<< obsm4 >>
rect -228 154 8 390
<< metal5 >>
rect 232 432 552 765
rect 872 432 1335 778
rect -252 112 552 432
rect 232 -221 552 112
rect 872 -234 1335 112
<< labels >>
rlabel locali s 28 215 248 255 6 A
port 1 nsew signal input
rlabel metal5 s 872 -234 1335 112 8 VGND
port 2 nsew ground bidirectional abutment
rlabel metal4 s 986 -179 1222 57 8 VGND
port 2 nsew ground bidirectional abutment
rlabel via3 s 1112 -32 1176 32 8 VGND
port 2 nsew ground bidirectional abutment
rlabel via3 s 1032 -32 1096 32 8 VGND
port 2 nsew ground bidirectional abutment
rlabel metal3 s 1026 -33 1182 33 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 1027 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 4 nsew power bidirectional
rlabel metal5 s 872 432 1335 778 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal4 s 986 487 1222 723 6 VPWR
port 5 nsew power bidirectional abutment
rlabel via3 s 1112 512 1176 576 6 VPWR
port 5 nsew power bidirectional abutment
rlabel via3 s 1032 512 1096 576 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal3 s 1026 511 1182 577 6 VPWR
port 5 nsew power bidirectional abutment
rlabel metal5 s 232 -221 552 112 8 X
port 6 nsew signal output
rlabel metal5 s -252 112 552 432 6 X
port 6 nsew signal output
rlabel metal5 s 232 432 552 765 6 X
port 6 nsew signal output
rlabel metal4 s 292 154 528 390 6 X
port 6 nsew signal output
rlabel via3 s 463 206 527 270 6 X
port 6 nsew signal output
rlabel via3 s 383 206 447 270 6 X
port 6 nsew signal output
rlabel metal3 s 377 205 533 271 6 X
port 6 nsew signal output
rlabel via2 s 467 210 523 266 6 X
port 6 nsew signal output
rlabel via2 s 387 210 443 266 6 X
port 6 nsew signal output
rlabel metal2 s 378 210 532 266 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1104 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 31774
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 18966
<< end >>
