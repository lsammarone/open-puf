magic
tech sky130B
magscale 1 2
timestamp 1648127584
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 732 203
rect 30 -17 64 21
<< scnmos >>
rect 80 47 110 177
rect 152 47 182 177
rect 339 47 369 177
rect 425 47 455 177
rect 519 47 549 177
rect 605 47 635 177
<< scpmoshvt >>
rect 80 297 110 497
rect 166 297 196 497
rect 343 297 373 497
rect 415 297 445 497
rect 523 297 553 497
rect 609 297 639 497
<< ndiff >>
rect 27 161 80 177
rect 27 127 36 161
rect 70 127 80 161
rect 27 93 80 127
rect 27 59 36 93
rect 70 59 80 93
rect 27 47 80 59
rect 110 47 152 177
rect 182 165 234 177
rect 182 131 192 165
rect 226 131 234 165
rect 182 120 234 131
rect 182 47 232 120
rect 289 104 339 177
rect 287 93 339 104
rect 287 59 295 93
rect 329 59 339 93
rect 287 47 339 59
rect 369 163 425 177
rect 369 129 380 163
rect 414 129 425 163
rect 369 47 425 129
rect 455 89 519 177
rect 455 55 470 89
rect 504 55 519 89
rect 455 47 519 55
rect 549 157 605 177
rect 549 123 560 157
rect 594 123 605 157
rect 549 89 605 123
rect 549 55 560 89
rect 594 55 605 89
rect 549 47 605 55
rect 635 89 706 177
rect 635 55 660 89
rect 694 55 706 89
rect 635 47 706 55
<< pdiff >>
rect 27 477 80 497
rect 27 443 35 477
rect 69 443 80 477
rect 27 381 80 443
rect 27 347 35 381
rect 69 347 80 381
rect 27 297 80 347
rect 110 489 166 497
rect 110 455 121 489
rect 155 455 166 489
rect 110 421 166 455
rect 110 387 121 421
rect 155 387 166 421
rect 110 297 166 387
rect 196 464 343 497
rect 196 430 221 464
rect 255 430 289 464
rect 323 430 343 464
rect 196 395 343 430
rect 196 361 221 395
rect 255 361 289 395
rect 323 361 343 395
rect 196 297 343 361
rect 373 297 415 497
rect 445 489 523 497
rect 445 455 466 489
rect 500 455 523 489
rect 445 421 523 455
rect 445 387 466 421
rect 500 387 523 421
rect 445 297 523 387
rect 553 477 609 497
rect 553 443 564 477
rect 598 443 609 477
rect 553 297 609 443
rect 639 485 692 497
rect 639 451 650 485
rect 684 451 692 485
rect 639 297 692 451
<< ndiffc >>
rect 36 127 70 161
rect 36 59 70 93
rect 192 131 226 165
rect 295 59 329 93
rect 380 129 414 163
rect 470 55 504 89
rect 560 123 594 157
rect 560 55 594 89
rect 660 55 694 89
<< pdiffc >>
rect 35 443 69 477
rect 35 347 69 381
rect 121 455 155 489
rect 121 387 155 421
rect 221 430 255 464
rect 289 430 323 464
rect 221 361 255 395
rect 289 361 323 395
rect 466 455 500 489
rect 466 387 500 421
rect 564 443 598 477
rect 650 451 684 485
<< poly >>
rect 80 497 110 523
rect 166 497 196 523
rect 343 497 373 523
rect 415 497 445 523
rect 523 497 553 523
rect 609 497 639 523
rect 80 274 110 297
rect 21 249 110 274
rect 166 265 196 297
rect 343 277 373 297
rect 21 215 38 249
rect 72 215 110 249
rect 21 199 110 215
rect 80 177 110 199
rect 152 249 220 265
rect 152 215 176 249
rect 210 215 220 249
rect 152 199 220 215
rect 295 249 373 277
rect 295 215 320 249
rect 354 215 373 249
rect 295 199 373 215
rect 415 265 445 297
rect 415 249 477 265
rect 523 264 553 297
rect 609 264 639 297
rect 415 215 431 249
rect 465 215 477 249
rect 415 199 477 215
rect 519 249 685 264
rect 519 215 533 249
rect 567 215 601 249
rect 635 215 685 249
rect 519 199 685 215
rect 152 177 182 199
rect 339 177 369 199
rect 425 177 455 199
rect 519 177 549 199
rect 605 177 635 199
rect 80 21 110 47
rect 152 21 182 47
rect 339 21 369 47
rect 425 21 455 47
rect 519 21 549 47
rect 605 21 635 47
<< polycont >>
rect 38 215 72 249
rect 176 215 210 249
rect 320 215 354 249
rect 431 215 465 249
rect 533 215 567 249
rect 601 215 635 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 18 477 71 493
rect 18 443 35 477
rect 69 443 71 477
rect 18 381 71 443
rect 105 489 171 527
rect 105 455 121 489
rect 155 455 171 489
rect 105 421 171 455
rect 105 387 121 421
rect 155 387 171 421
rect 205 464 339 493
rect 205 430 221 464
rect 255 430 289 464
rect 323 430 339 464
rect 205 395 339 430
rect 18 347 35 381
rect 69 353 71 381
rect 205 361 221 395
rect 255 361 289 395
rect 323 361 339 395
rect 440 489 526 527
rect 440 455 466 489
rect 500 455 526 489
rect 440 421 526 455
rect 440 387 466 421
rect 500 387 526 421
rect 562 477 600 493
rect 562 443 564 477
rect 598 443 600 477
rect 634 485 700 527
rect 634 451 650 485
rect 684 451 700 485
rect 562 415 600 443
rect 562 381 708 415
rect 205 353 339 361
rect 69 347 533 353
rect 18 302 533 347
rect 17 249 72 265
rect 17 215 38 249
rect 17 199 72 215
rect 106 165 142 302
rect 499 265 533 302
rect 176 249 248 265
rect 210 215 248 249
rect 176 199 248 215
rect 306 249 364 265
rect 306 215 320 249
rect 354 215 364 249
rect 306 199 364 215
rect 398 249 465 265
rect 398 215 431 249
rect 398 199 465 215
rect 499 249 635 265
rect 499 215 533 249
rect 567 215 601 249
rect 499 199 635 215
rect 19 161 142 165
rect 19 127 36 161
rect 70 127 142 161
rect 176 131 192 165
rect 226 163 430 165
rect 226 131 380 163
rect 176 129 380 131
rect 414 129 430 163
rect 669 157 708 381
rect 176 127 430 129
rect 19 93 142 127
rect 544 123 560 157
rect 594 123 708 157
rect 19 59 36 93
rect 70 85 142 93
rect 70 59 86 85
rect 19 51 86 59
rect 278 59 295 93
rect 329 59 345 93
rect 278 17 345 59
rect 463 89 510 105
rect 463 55 470 89
rect 504 55 510 89
rect 463 17 510 55
rect 544 89 610 123
rect 544 55 560 89
rect 594 55 610 89
rect 544 51 610 55
rect 644 55 660 89
rect 694 55 710 89
rect 644 17 710 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 674 153 708 187 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 o211a_2
rlabel metal1 s 0 -48 736 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 770980
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 764656
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 3.680 0.000 
<< end >>
