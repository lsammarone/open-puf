/farmshare/home/classes/ee/372/PDKs/share/pdk/sky130A/libs.tech/ngspice/sky130_fd_pr__model__diode_pd2nw_11v0.model.spice