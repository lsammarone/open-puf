/farmshare/home/classes/ee/372/PDKs/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_01v8.pm3.spice